
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

use work.ctp7_utils_pkg.all;


library UNISIM;
use UNISIM.VCOMPONENTS.all;

entity ctp7_top is
  generic (
    C_DATE_CODE      : std_logic_vector (31 downto 0) := x"00000000";
    C_GITHASH_CODE   : std_logic_vector (31 downto 0) := x"00000000";
    C_GIT_REPO_DIRTY : std_logic                      := '0'
    );
  Port (
  
      clk_200_diff_in_clk_p : in std_logic;
      clk_200_diff_in_clk_n : in std_logic;
    
      LEDs : out std_logic_vector (1 downto 0);
    
      LED_GREEN_o : out std_logic;
      LED_RED_o   : out std_logic;
      LED_BLUE_o  : out std_logic;
    
      axi_c2c_v7_to_zynq_data        : out std_logic_vector (16 downto 0);
      axi_c2c_v7_to_zynq_clk         : out std_logic;
      axi_c2c_zynq_to_v7_clk         : in  std_logic;
      axi_c2c_zynq_to_v7_data        : in  std_logic_vector (16 downto 0);
      axi_c2c_v7_to_zynq_link_status : out std_logic;
      axi_c2c_zynq_to_v7_reset       : in  std_logic
   );
end ctp7_top;

architecture ctp7_top_arch of ctp7_top is

  component v7_bd is
  port (

    clk_200_diff_in_clk_n : in STD_LOGIC;
    clk_200_diff_in_clk_p : in STD_LOGIC;
    
    axi_c2c_zynq_to_v7_clk : in STD_LOGIC;
    axi_c2c_zynq_to_v7_data : in STD_LOGIC_VECTOR ( 16 downto 0 );
    axi_c2c_v7_to_zynq_link_status : out STD_LOGIC;
    axi_c2c_v7_to_zynq_clk : out STD_LOGIC;
    axi_c2c_v7_to_zynq_data : out STD_LOGIC_VECTOR ( 16 downto 0 );
    axi_c2c_zynq_to_v7_reset : in STD_LOGIC;

    BRAM_CTRL_REG_FILE_addr : out STD_LOGIC_VECTOR ( 16 downto 0 );
    BRAM_CTRL_REG_FILE_clk : out STD_LOGIC;
    BRAM_CTRL_REG_FILE_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_REG_FILE_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_REG_FILE_en : out STD_LOGIC;
    BRAM_CTRL_REG_FILE_rst : out STD_LOGIC;
    BRAM_CTRL_REG_FILE_we : out STD_LOGIC_VECTOR ( 3 downto 0 );

    BRAM_CTRL_INPUT_RAM_0_addr : out STD_LOGIC_VECTOR ( 16 downto 0 );
    BRAM_CTRL_INPUT_RAM_0_clk : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_0_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_INPUT_RAM_0_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_INPUT_RAM_0_en : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_0_rst : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_0_we : out STD_LOGIC_VECTOR ( 3 downto 0 );

    BRAM_CTRL_INPUT_RAM_1_addr : out STD_LOGIC_VECTOR ( 16 downto 0 );
    BRAM_CTRL_INPUT_RAM_1_clk : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_1_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_INPUT_RAM_1_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_INPUT_RAM_1_en : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_1_rst : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_1_we : out STD_LOGIC_VECTOR ( 3 downto 0 );
    
    BRAM_CTRL_INPUT_RAM_2_addr : out STD_LOGIC_VECTOR ( 16 downto 0 );
    BRAM_CTRL_INPUT_RAM_2_clk : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_2_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_INPUT_RAM_2_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_INPUT_RAM_2_en : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_2_rst : out STD_LOGIC;
    BRAM_CTRL_INPUT_RAM_2_we : out STD_LOGIC_VECTOR ( 3 downto 0 );
    
    BRAM_CTRL_OUTPUT_RAM_0_addr : out STD_LOGIC_VECTOR ( 16 downto 0 );
    BRAM_CTRL_OUTPUT_RAM_0_clk : out STD_LOGIC;
    BRAM_CTRL_OUTPUT_RAM_0_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_OUTPUT_RAM_0_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_OUTPUT_RAM_0_en : out STD_LOGIC;
    BRAM_CTRL_OUTPUT_RAM_0_rst : out STD_LOGIC;
    BRAM_CTRL_OUTPUT_RAM_0_we : out STD_LOGIC_VECTOR ( 3 downto 0 );
    
    BRAM_CTRL_OUTPUT_RAM_1_addr : out STD_LOGIC_VECTOR ( 16 downto 0 );
    BRAM_CTRL_OUTPUT_RAM_1_clk : out STD_LOGIC;
    BRAM_CTRL_OUTPUT_RAM_1_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_OUTPUT_RAM_1_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    BRAM_CTRL_OUTPUT_RAM_1_en : out STD_LOGIC;
    BRAM_CTRL_OUTPUT_RAM_1_rst : out STD_LOGIC;
    BRAM_CTRL_OUTPUT_RAM_1_we : out STD_LOGIC_VECTOR ( 3 downto 0 );
    
    clk_50mhz : out STD_LOGIC;
    clk_240mhz : out STD_LOGIC    
    
  );
  end component v7_bd;
  
COMPONENT ila_hls
       
       PORT (
           clk : IN STD_LOGIC;
       
       
       
           probe0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
           probe1 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
           probe2 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
           probe3 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
           probe4 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
           probe5 : IN STD_LOGIC_VECTOR(0 DOWNTO 0); 
           probe6 : IN STD_LOGIC_VECTOR(191 DOWNTO 0);
           probe7 : IN STD_LOGIC_VECTOR(191 DOWNTO 0)
       );
       END COMPONENT  ;
  

  signal s_clk_50  : std_logic;
  signal s_clk_240        : std_logic;

  signal BRAM_CTRL_REG_FILE_en   : std_logic;
  signal BRAM_CTRL_REG_FILE_dout : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_REG_FILE_din  : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_REG_FILE_we   : std_logic_vector (3 downto 0);
  signal BRAM_CTRL_REG_FILE_addr : std_logic_vector (16 downto 0);
  signal BRAM_CTRL_REG_FILE_clk  : std_logic;
  signal BRAM_CTRL_REG_FILE_rst  : std_logic;

  signal BRAM_CTRL_INPUT_RAM_0_addr : std_logic_vector (16 downto 0);
  signal BRAM_CTRL_INPUT_RAM_0_clk  : std_logic;
  signal BRAM_CTRL_INPUT_RAM_0_din  : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_INPUT_RAM_0_dout : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_INPUT_RAM_0_en   : std_logic;
  signal BRAM_CTRL_INPUT_RAM_0_rst  : std_logic;
  signal BRAM_CTRL_INPUT_RAM_0_we   : std_logic_vector (3 downto 0);

  signal BRAM_CTRL_INPUT_RAM_1_addr : std_logic_vector (16 downto 0);
  signal BRAM_CTRL_INPUT_RAM_1_clk  : std_logic;
  signal BRAM_CTRL_INPUT_RAM_1_din  : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_INPUT_RAM_1_dout : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_INPUT_RAM_1_en   : std_logic;
  signal BRAM_CTRL_INPUT_RAM_1_rst  : std_logic;
  signal BRAM_CTRL_INPUT_RAM_1_we   : std_logic_vector (3 downto 0);
  
  signal BRAM_CTRL_INPUT_RAM_2_addr : std_logic_vector (16 downto 0);
  signal BRAM_CTRL_INPUT_RAM_2_clk  : std_logic;
  signal BRAM_CTRL_INPUT_RAM_2_din  : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_INPUT_RAM_2_dout : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_INPUT_RAM_2_en   : std_logic;
  signal BRAM_CTRL_INPUT_RAM_2_rst  : std_logic;
  signal BRAM_CTRL_INPUT_RAM_2_we   : std_logic_vector (3 downto 0);

  signal BRAM_CTRL_OUTPUT_RAM_0_addr : std_logic_vector (16 downto 0); 
  signal BRAM_CTRL_OUTPUT_RAM_0_clk  : std_logic;
  signal BRAM_CTRL_OUTPUT_RAM_0_din  : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_OUTPUT_RAM_0_dout : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_OUTPUT_RAM_0_en   : std_logic;
  signal BRAM_CTRL_OUTPUT_RAM_0_rst  : std_logic;
  signal BRAM_CTRL_OUTPUT_RAM_0_we   : std_logic_vector (3 downto 0);

  signal BRAM_CTRL_OUTPUT_RAM_1_addr : std_logic_vector (16 downto 0);
  signal BRAM_CTRL_OUTPUT_RAM_1_clk  : std_logic;
  signal BRAM_CTRL_OUTPUT_RAM_1_din  : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_OUTPUT_RAM_1_dout : std_logic_vector (31 downto 0);
  signal BRAM_CTRL_OUTPUT_RAM_1_en   : std_logic;
  signal BRAM_CTRL_OUTPUT_RAM_1_rst  : std_logic;
  signal BRAM_CTRL_OUTPUT_RAM_1_we   : std_logic_vector (3 downto 0);

  signal s_LED_FP : std_logic_vector(31 downto 0);
  
  signal s_pattern_start_request: std_logic;
  signal s_algo_latency :  std_logic_vector ( 15 downto 0 );
  
  signal s_pattern_start, s_pattern_start_s1, s_pattern_start_s2:  std_logic;
  
  signal s_INPUT_RAM_start:  std_logic;
  signal s_OUTPUT_RAM_start:  std_logic;
  
  signal s_INPUT_link_arr :  t_slv_arr_192(66 downto 0) := (others => (others => '0'));
  signal s_OUTPUT_link_arr:   t_slv_arr_192(47 downto 0) := (others => (others => '0'));
  signal s_cfg_reg : t_slv_arr_32(31 downto 0);

-----------------------------------------------------------------------------
-- Begin User_Code
-----------------------------------------------------------------------------
 COMPONENT Getclustertracklinker_3
    PORT (
      ap_clk : IN STD_LOGIC;
      ap_rst : IN STD_LOGIC;
      ap_start : IN STD_LOGIC;
      ap_done : OUT STD_LOGIC;
      ap_idle : OUT STD_LOGIC;
      ap_ready : OUT STD_LOGIC;
      
      ClusterET_0_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_0_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_0_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_0_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_1_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_1_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_1_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_1_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_2_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_2_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_2_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_2_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_3_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_3_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_3_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_3_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_4_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_4_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_4_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_4_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_5_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_5_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_5_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_5_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_6_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_6_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_6_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_6_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_7_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_7_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_7_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_7_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_8_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_8_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_8_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_8_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_9_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_9_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_9_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_9_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_10_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_10_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_10_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_10_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_11_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_11_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_11_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_11_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_12_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_12_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_12_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_12_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_13_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_13_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_13_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_13_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_14_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_14_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_14_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_14_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_15_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_15_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_15_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_15_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_16_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_16_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_16_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      ClusterET_16_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      
      
      peakEta_0_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_0_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_0_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_0_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_1_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_1_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_1_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_1_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_2_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_2_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_2_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_2_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_3_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_3_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_3_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_3_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_4_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_4_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_4_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_4_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_5_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_5_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_5_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_5_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_6_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_6_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_6_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_6_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_7_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_7_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_7_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_7_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_8_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_8_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_8_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_8_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_9_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_9_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_9_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_9_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_10_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_10_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_10_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_10_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_11_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_11_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_11_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_11_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_12_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_12_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_12_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_12_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_13_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_13_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_13_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_13_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_14_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_14_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_14_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_14_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_15_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_15_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_15_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_15_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_16_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_16_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_16_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakEta_16_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      
      
      peakPhi_0_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_0_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_0_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_0_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_1_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_1_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_1_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_1_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_2_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_2_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_2_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_2_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_3_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_3_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_3_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_3_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_4_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_4_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_4_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_4_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_5_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_5_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_5_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_5_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_6_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_6_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_6_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_6_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_7_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_7_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_7_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_7_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_8_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_8_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_8_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_8_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_9_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_9_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_9_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_9_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_10_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_10_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_10_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_10_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_11_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_11_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_11_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_11_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_12_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_12_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_12_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_12_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_13_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_13_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_13_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_13_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_14_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_14_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_14_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_14_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_15_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_15_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_15_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_15_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_16_0_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_16_1_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_16_2_V : IN STD_LOGIC_VECTOR (2 downto 0);
      peakPhi_16_3_V : IN STD_LOGIC_VECTOR (2 downto 0);
      
      
      trackPT_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_4_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_5_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_6_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_7_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_8_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPT_9_V : IN STD_LOGIC_VECTOR (9 downto 0);
      
      
      trackEta_0_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_1_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_2_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_3_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_4_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_5_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_6_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_7_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_8_V : IN STD_LOGIC_VECTOR (8 downto 0);
      trackEta_9_V : IN STD_LOGIC_VECTOR (8 downto 0);
      
      
      trackPhi_0_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_1_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_2_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_3_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_4_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_5_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_6_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_7_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_8_V : IN STD_LOGIC_VECTOR (9 downto 0);
      trackPhi_9_V : IN STD_LOGIC_VECTOR (9 downto 0);
      
      
      output_linkedTrackPT_0_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_1_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_2_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_3_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_4_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_5_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_6_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_7_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_8_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPT_9_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      
      
      output_linkedTrackEta_0_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_1_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_2_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_3_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_4_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_5_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_6_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_7_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_8_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_linkedTrackEta_9_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      
      
      output_linkedTrackPhi_0_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_1_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_2_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_3_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_4_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_5_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_6_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_7_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_8_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_linkedTrackPhi_9_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      
      
      output_linkedTrackQuality_0_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_1_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_2_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_3_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_4_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_5_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_6_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_7_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_8_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      output_linkedTrackQuality_9_V : OUT STD_LOGIC_VECTOR (7 downto 0);
      
      
      output_neutralClusterET_0_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_1_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_2_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_3_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_4_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_5_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_6_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_7_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_8_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_9_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_10_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_11_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_12_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_13_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_14_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_15_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_16_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_17_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_18_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_19_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_20_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_21_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_22_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_23_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_24_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_25_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_26_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_27_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_28_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_29_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_30_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_31_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_32_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_33_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_34_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_35_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_36_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_37_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_38_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_39_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_40_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_41_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_42_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_43_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_44_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_45_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_46_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_47_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_48_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_49_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_50_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_51_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_52_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_53_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_54_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_55_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_56_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_57_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_58_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_59_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_60_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_61_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_62_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_63_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_64_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_65_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_66_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterET_67_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      
      
      output_neutralClusterEta_0_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_1_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_2_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_3_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_4_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_5_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_6_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_7_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_8_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_9_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_10_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_11_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_12_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_13_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_14_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_15_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_16_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_17_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_18_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_19_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_20_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_21_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_22_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_23_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_24_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_25_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_26_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_27_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_28_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_29_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_30_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_31_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_32_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_33_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_34_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_35_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_36_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_37_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_38_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_39_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_40_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_41_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_42_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_43_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_44_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_45_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_46_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_47_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_48_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_49_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_50_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_51_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_52_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_53_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_54_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_55_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_56_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_57_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_58_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_59_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_60_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_61_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_62_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_63_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_64_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_65_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_66_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      output_neutralClusterEta_67_V : OUT STD_LOGIC_VECTOR (8 downto 0);
      
      
      output_neutralClusterPhi_0_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_1_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_2_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_3_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_4_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_5_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_6_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_7_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_8_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_9_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_10_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_11_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_12_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_13_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_14_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_15_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_16_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_17_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_18_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_19_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_20_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_21_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_22_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_23_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_24_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_25_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_26_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_27_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_28_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_29_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_30_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_31_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_32_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_33_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_34_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_35_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_36_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_37_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_38_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_39_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_40_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_41_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_42_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_43_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_44_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_45_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_46_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_47_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_48_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_49_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_50_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_51_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_52_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_53_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_54_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_55_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_56_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_57_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_58_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_59_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_60_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_61_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_62_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_63_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_64_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_65_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_66_V : OUT STD_LOGIC_VECTOR (9 downto 0);
      output_neutralClusterPhi_67_V : OUT STD_LOGIC_VECTOR (9 downto 0)
    );
  END COMPONENT;  

-- HLS Algo Control/Handshake Interface
      signal ap_clk :  STD_LOGIC;
      signal ap_rst :  STD_LOGIC;
      signal ap_start :  STD_LOGIC;
      signal ap_done :  STD_LOGIC;
      signal ap_idle :  STD_LOGIC;
      signal ap_ready :  STD_LOGIC;
      
     
     signal ClusterET_0_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_0_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_0_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_0_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_1_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_1_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_1_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_1_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_2_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_2_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_2_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_2_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_3_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_3_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_3_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_3_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_4_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_4_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_4_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_4_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_5_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_5_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_5_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_5_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_6_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_6_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_6_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_6_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_7_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_7_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_7_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_7_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_8_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_8_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_8_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_8_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_9_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_9_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_9_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_9_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_10_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_10_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_10_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_10_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_11_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_11_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_11_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_11_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_12_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_12_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_12_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_12_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_13_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_13_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_13_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_13_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_14_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_14_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_14_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_14_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_15_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_15_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_15_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_15_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_16_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_16_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_16_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal ClusterET_16_3_V : STD_LOGIC_VECTOR (9 downto 0);
      
      
      signal peakEta_0_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_0_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_0_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_0_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_1_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_1_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_1_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_1_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_2_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_2_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_2_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_2_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_3_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_3_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_3_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_3_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_4_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_4_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_4_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_4_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_5_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_5_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_5_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_5_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_6_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_6_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_6_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_6_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_7_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_7_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_7_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_7_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_8_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_8_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_8_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_8_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_9_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_9_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_9_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_9_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_10_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_10_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_10_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_10_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_11_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_11_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_11_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_11_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_12_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_12_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_12_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_12_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_13_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_13_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_13_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_13_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_14_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_14_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_14_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_14_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_15_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_15_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_15_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_15_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_16_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_16_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_16_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakEta_16_3_V : STD_LOGIC_VECTOR (2 downto 0);
      
      
      signal peakPhi_0_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_0_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_0_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_0_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_1_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_1_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_1_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_1_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_2_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_2_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_2_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_2_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_3_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_3_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_3_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_3_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_4_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_4_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_4_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_4_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_5_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_5_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_5_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_5_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_6_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_6_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_6_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_6_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_7_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_7_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_7_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_7_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_8_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_8_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_8_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_8_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_9_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_9_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_9_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_9_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_10_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_10_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_10_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_10_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_11_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_11_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_11_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_11_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_12_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_12_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_12_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_12_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_13_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_13_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_13_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_13_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_14_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_14_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_14_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_14_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_15_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_15_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_15_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_15_3_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_16_0_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_16_1_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_16_2_V : STD_LOGIC_VECTOR (2 downto 0);
      signal peakPhi_16_3_V : STD_LOGIC_VECTOR (2 downto 0);
      
      
      signal trackPT_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_4_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_5_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_6_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_7_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_8_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPT_9_V : STD_LOGIC_VECTOR (9 downto 0);
      
      
      signal trackEta_0_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_1_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_2_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_3_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_4_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_5_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_6_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_7_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_8_V : STD_LOGIC_VECTOR (8 downto 0);
      signal trackEta_9_V : STD_LOGIC_VECTOR (8 downto 0);
      
      
      signal trackPhi_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_4_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_5_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_6_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_7_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_8_V : STD_LOGIC_VECTOR (9 downto 0);
      signal trackPhi_9_V : STD_LOGIC_VECTOR (9 downto 0);
      
      
      signal output_linkedTrackPT_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_4_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_5_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_6_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_7_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_8_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPT_9_V : STD_LOGIC_VECTOR (9 downto 0);
      
      
      signal output_linkedTrackEta_0_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_1_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_2_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_3_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_4_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_5_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_6_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_7_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_8_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_linkedTrackEta_9_V : STD_LOGIC_VECTOR (8 downto 0);
      
      
      signal output_linkedTrackPhi_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_4_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_5_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_6_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_7_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_8_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_linkedTrackPhi_9_V : STD_LOGIC_VECTOR (9 downto 0);
      
      
      signal output_linkedTrackQuality_0_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_1_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_2_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_3_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_4_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_5_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_6_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_7_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_8_V : STD_LOGIC_VECTOR (7 downto 0);
      signal output_linkedTrackQuality_9_V : STD_LOGIC_VECTOR (7 downto 0);
      
      
      signal output_neutralClusterET_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_4_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_5_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_6_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_7_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_8_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_9_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_10_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_11_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_12_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_13_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_14_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_15_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_16_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_17_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_18_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_19_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_20_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_21_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_22_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_23_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_24_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_25_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_26_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_27_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_28_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_29_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_30_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_31_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_32_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_33_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_34_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_35_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_36_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_37_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_38_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_39_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_40_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_41_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_42_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_43_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_44_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_45_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_46_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_47_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_48_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_49_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_50_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_51_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_52_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_53_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_54_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_55_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_56_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_57_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_58_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_59_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_60_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_61_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_62_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_63_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_64_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_65_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_66_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterET_67_V : STD_LOGIC_VECTOR (9 downto 0);
      
      
      signal output_neutralClusterEta_0_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_1_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_2_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_3_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_4_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_5_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_6_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_7_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_8_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_9_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_10_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_11_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_12_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_13_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_14_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_15_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_16_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_17_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_18_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_19_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_20_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_21_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_22_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_23_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_24_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_25_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_26_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_27_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_28_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_29_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_30_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_31_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_32_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_33_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_34_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_35_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_36_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_37_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_38_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_39_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_40_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_41_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_42_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_43_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_44_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_45_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_46_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_47_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_48_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_49_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_50_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_51_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_52_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_53_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_54_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_55_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_56_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_57_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_58_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_59_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_60_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_61_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_62_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_63_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_64_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_65_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_66_V : STD_LOGIC_VECTOR (8 downto 0);
      signal output_neutralClusterEta_67_V : STD_LOGIC_VECTOR (8 downto 0);
      
      
      signal output_neutralClusterPhi_0_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_1_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_2_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_3_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_4_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_5_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_6_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_7_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_8_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_9_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_10_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_11_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_12_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_13_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_14_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_15_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_16_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_17_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_18_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_19_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_20_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_21_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_22_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_23_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_24_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_25_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_26_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_27_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_28_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_29_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_30_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_31_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_32_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_33_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_34_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_35_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_36_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_37_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_38_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_39_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_40_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_41_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_42_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_43_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_44_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_45_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_46_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_47_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_48_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_49_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_50_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_51_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_52_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_53_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_54_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_55_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_56_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_57_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_58_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_59_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_60_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_61_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_62_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_63_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_64_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_65_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_66_V : STD_LOGIC_VECTOR (9 downto 0);
      signal output_neutralClusterPhi_67_V : STD_LOGIC_VECTOR (9 downto 0);
      
-----------------------------------------------------------------------------
-- End User_Code
-----------------------------------------------------------------------------
           
begin

    LED_GREEN_o <= s_LED_FP(0);
    LED_RED_o   <= s_LED_FP(1);
    LED_BLUE_o  <= s_LED_FP(2);

  i_v7_bd : v7_bd
    port map (
    
        axi_c2c_v7_to_zynq_clk               => axi_c2c_v7_to_zynq_clk,
        axi_c2c_v7_to_zynq_data(16 downto 0) => axi_c2c_v7_to_zynq_data(16 downto 0),
        axi_c2c_v7_to_zynq_link_status       => axi_c2c_v7_to_zynq_link_status,
        axi_c2c_zynq_to_v7_clk               => axi_c2c_zynq_to_v7_clk,
        axi_c2c_zynq_to_v7_data(16 downto 0) => axi_c2c_zynq_to_v7_data(16 downto 0),
        axi_c2c_zynq_to_v7_reset             => axi_c2c_zynq_to_v7_reset,
    
        clk_200_diff_in_clk_n => clk_200_diff_in_clk_n,
        clk_200_diff_in_clk_p => clk_200_diff_in_clk_p,
        
        BRAM_CTRL_REG_FILE_addr => BRAM_CTRL_REG_FILE_addr,
        BRAM_CTRL_REG_FILE_clk  => BRAM_CTRL_REG_FILE_clk,
        BRAM_CTRL_REG_FILE_din  => BRAM_CTRL_REG_FILE_din,
        BRAM_CTRL_REG_FILE_dout => BRAM_CTRL_REG_FILE_dout,
        BRAM_CTRL_REG_FILE_en   => BRAM_CTRL_REG_FILE_en,
        BRAM_CTRL_REG_FILE_rst  => BRAM_CTRL_REG_FILE_rst,
        BRAM_CTRL_REG_FILE_we   => BRAM_CTRL_REG_FILE_we,

        BRAM_CTRL_INPUT_RAM_0_addr => BRAM_CTRL_INPUT_RAM_0_addr,
        BRAM_CTRL_INPUT_RAM_0_clk  => BRAM_CTRL_INPUT_RAM_0_clk,
        BRAM_CTRL_INPUT_RAM_0_din  => BRAM_CTRL_INPUT_RAM_0_din,
        BRAM_CTRL_INPUT_RAM_0_dout => BRAM_CTRL_INPUT_RAM_0_dout,
        BRAM_CTRL_INPUT_RAM_0_en   => BRAM_CTRL_INPUT_RAM_0_en,
        BRAM_CTRL_INPUT_RAM_0_rst  => BRAM_CTRL_INPUT_RAM_0_rst,
        BRAM_CTRL_INPUT_RAM_0_we   => BRAM_CTRL_INPUT_RAM_0_we,

        BRAM_CTRL_INPUT_RAM_1_addr => BRAM_CTRL_INPUT_RAM_1_addr,
        BRAM_CTRL_INPUT_RAM_1_clk  => BRAM_CTRL_INPUT_RAM_1_clk,
        BRAM_CTRL_INPUT_RAM_1_din  => BRAM_CTRL_INPUT_RAM_1_din,
        BRAM_CTRL_INPUT_RAM_1_dout => BRAM_CTRL_INPUT_RAM_1_dout,
        BRAM_CTRL_INPUT_RAM_1_en   => BRAM_CTRL_INPUT_RAM_1_en,
        BRAM_CTRL_INPUT_RAM_1_rst  => BRAM_CTRL_INPUT_RAM_1_rst,
        BRAM_CTRL_INPUT_RAM_1_we   => BRAM_CTRL_INPUT_RAM_1_we,
        
        BRAM_CTRL_INPUT_RAM_2_addr => BRAM_CTRL_INPUT_RAM_2_addr,
        BRAM_CTRL_INPUT_RAM_2_clk  => BRAM_CTRL_INPUT_RAM_2_clk,
        BRAM_CTRL_INPUT_RAM_2_din  => BRAM_CTRL_INPUT_RAM_2_din,
        BRAM_CTRL_INPUT_RAM_2_dout => BRAM_CTRL_INPUT_RAM_2_dout,
        BRAM_CTRL_INPUT_RAM_2_en   => BRAM_CTRL_INPUT_RAM_2_en,
        BRAM_CTRL_INPUT_RAM_2_rst  => BRAM_CTRL_INPUT_RAM_2_rst,
        BRAM_CTRL_INPUT_RAM_2_we   => BRAM_CTRL_INPUT_RAM_2_we,
        
        BRAM_CTRL_OUTPUT_RAM_0_addr => BRAM_CTRL_OUTPUT_RAM_0_addr,
        BRAM_CTRL_OUTPUT_RAM_0_clk  => BRAM_CTRL_OUTPUT_RAM_0_clk,
        BRAM_CTRL_OUTPUT_RAM_0_din  => BRAM_CTRL_OUTPUT_RAM_0_din,
        BRAM_CTRL_OUTPUT_RAM_0_dout => BRAM_CTRL_OUTPUT_RAM_0_dout,
        BRAM_CTRL_OUTPUT_RAM_0_en   => BRAM_CTRL_OUTPUT_RAM_0_en,
        BRAM_CTRL_OUTPUT_RAM_0_rst  => BRAM_CTRL_OUTPUT_RAM_0_rst,
        BRAM_CTRL_OUTPUT_RAM_0_we   => BRAM_CTRL_OUTPUT_RAM_0_we,
 
        BRAM_CTRL_OUTPUT_RAM_1_addr => BRAM_CTRL_OUTPUT_RAM_1_addr,
        BRAM_CTRL_OUTPUT_RAM_1_clk  => BRAM_CTRL_OUTPUT_RAM_1_clk,
        BRAM_CTRL_OUTPUT_RAM_1_din  => BRAM_CTRL_OUTPUT_RAM_1_din,
        BRAM_CTRL_OUTPUT_RAM_1_dout => BRAM_CTRL_OUTPUT_RAM_1_dout,
        BRAM_CTRL_OUTPUT_RAM_1_en   => BRAM_CTRL_OUTPUT_RAM_1_en,
        BRAM_CTRL_OUTPUT_RAM_1_rst  => BRAM_CTRL_OUTPUT_RAM_1_rst,
        BRAM_CTRL_OUTPUT_RAM_1_we   => BRAM_CTRL_OUTPUT_RAM_1_we,        
        
        clk_50mhz  => s_clk_50,
        clk_240mhz => s_clk_240
      );
      
  i_register_file : entity work.register_file
        generic map(
          C_DATE_CODE      => C_DATE_CODE,
          C_GITHASH_CODE   => C_GITHASH_CODE,
          C_GIT_REPO_DIRTY => C_GIT_REPO_DIRTY
          )
        port map (
    
          LED_FP_o => s_led_FP,
   
          BRAM_CTRL_REG_FILE_addr => BRAM_CTRL_REG_FILE_addr,
          BRAM_CTRL_REG_FILE_clk  => BRAM_CTRL_REG_FILE_clk,
          BRAM_CTRL_REG_FILE_din  => BRAM_CTRL_REG_FILE_din,
          BRAM_CTRL_REG_FILE_dout => BRAM_CTRL_REG_FILE_dout,
          BRAM_CTRL_REG_FILE_en   => BRAM_CTRL_REG_FILE_en,
          BRAM_CTRL_REG_FILE_rst  => BRAM_CTRL_REG_FILE_rst,
          BRAM_CTRL_REG_FILE_we   => BRAM_CTRL_REG_FILE_we,
          
          pattern_start_o => s_pattern_start,
          cfg_reg_o  => s_cfg_reg

          );   
          
s_pattern_start_s1 <= s_pattern_start when rising_edge(s_clk_240);
s_pattern_start_s2 <= s_pattern_start_s1 when rising_edge(s_clk_240);

          
i_pattern_io_engine : entity work.pattern_io_engine 
    Port map( 
    
        clk_240_i => s_clk_240,
        
        pattern_restart_i  => s_pattern_start_s2,
        
        algo_rst_o  => ap_rst,
        algo_start_o  => ap_start,
        algo_done_i  => ap_done,
        
        INPUT_link_arr_o  => s_INPUT_link_arr,
        OUTPUT_link_arr_i => s_OUTPUT_link_arr,
        
        BRAM_CTRL_INPUT_RAM_0_addr => BRAM_CTRL_INPUT_RAM_0_addr,
        BRAM_CTRL_INPUT_RAM_0_clk  => BRAM_CTRL_INPUT_RAM_0_clk,
        BRAM_CTRL_INPUT_RAM_0_din  => BRAM_CTRL_INPUT_RAM_0_din,
        BRAM_CTRL_INPUT_RAM_0_dout => BRAM_CTRL_INPUT_RAM_0_dout,
        BRAM_CTRL_INPUT_RAM_0_en   => BRAM_CTRL_INPUT_RAM_0_en,
        BRAM_CTRL_INPUT_RAM_0_rst  => BRAM_CTRL_INPUT_RAM_0_rst,
        BRAM_CTRL_INPUT_RAM_0_we   => BRAM_CTRL_INPUT_RAM_0_we,

        BRAM_CTRL_INPUT_RAM_1_addr => BRAM_CTRL_INPUT_RAM_1_addr,
        BRAM_CTRL_INPUT_RAM_1_clk  => BRAM_CTRL_INPUT_RAM_1_clk,
        BRAM_CTRL_INPUT_RAM_1_din  => BRAM_CTRL_INPUT_RAM_1_din,
        BRAM_CTRL_INPUT_RAM_1_dout => BRAM_CTRL_INPUT_RAM_1_dout,
        BRAM_CTRL_INPUT_RAM_1_en   => BRAM_CTRL_INPUT_RAM_1_en,
        BRAM_CTRL_INPUT_RAM_1_rst  => BRAM_CTRL_INPUT_RAM_1_rst,
        BRAM_CTRL_INPUT_RAM_1_we   => BRAM_CTRL_INPUT_RAM_1_we,
        
        BRAM_CTRL_INPUT_RAM_2_addr => BRAM_CTRL_INPUT_RAM_2_addr,
        BRAM_CTRL_INPUT_RAM_2_clk  => BRAM_CTRL_INPUT_RAM_2_clk,
        BRAM_CTRL_INPUT_RAM_2_din  => BRAM_CTRL_INPUT_RAM_2_din,
        BRAM_CTRL_INPUT_RAM_2_dout => BRAM_CTRL_INPUT_RAM_2_dout,
        BRAM_CTRL_INPUT_RAM_2_en   => BRAM_CTRL_INPUT_RAM_2_en,
        BRAM_CTRL_INPUT_RAM_2_rst  => BRAM_CTRL_INPUT_RAM_2_rst,
        BRAM_CTRL_INPUT_RAM_2_we   => BRAM_CTRL_INPUT_RAM_2_we,
        
        BRAM_CTRL_OUTPUT_RAM_0_addr => BRAM_CTRL_OUTPUT_RAM_0_addr,
        BRAM_CTRL_OUTPUT_RAM_0_clk  => BRAM_CTRL_OUTPUT_RAM_0_clk,
        BRAM_CTRL_OUTPUT_RAM_0_din  => BRAM_CTRL_OUTPUT_RAM_0_din,
        BRAM_CTRL_OUTPUT_RAM_0_dout => BRAM_CTRL_OUTPUT_RAM_0_dout,
        BRAM_CTRL_OUTPUT_RAM_0_en   => BRAM_CTRL_OUTPUT_RAM_0_en,
        BRAM_CTRL_OUTPUT_RAM_0_rst  => BRAM_CTRL_OUTPUT_RAM_0_rst,
        BRAM_CTRL_OUTPUT_RAM_0_we   => BRAM_CTRL_OUTPUT_RAM_0_we,
 
        BRAM_CTRL_OUTPUT_RAM_1_addr => BRAM_CTRL_OUTPUT_RAM_1_addr,
        BRAM_CTRL_OUTPUT_RAM_1_clk  => BRAM_CTRL_OUTPUT_RAM_1_clk,
        BRAM_CTRL_OUTPUT_RAM_1_din  => BRAM_CTRL_OUTPUT_RAM_1_din,
        BRAM_CTRL_OUTPUT_RAM_1_dout => BRAM_CTRL_OUTPUT_RAM_1_dout,
        BRAM_CTRL_OUTPUT_RAM_1_en   => BRAM_CTRL_OUTPUT_RAM_1_en,
        BRAM_CTRL_OUTPUT_RAM_1_rst  => BRAM_CTRL_OUTPUT_RAM_1_rst,
        BRAM_CTRL_OUTPUT_RAM_1_we   => BRAM_CTRL_OUTPUT_RAM_1_we
     );          
     
     ap_clk <= s_clk_240; 
     
     i_ila_hls : ila_hls
     PORT MAP (
         clk => s_clk_240,     
         probe0(0) => ap_rst, 
         probe1(0) => ap_rst, 
         probe2(0) => ap_start, 
         probe3(0) => ap_done, 
         probe4(0) => ap_idle, 
         probe5(0) => ap_ready, 
         probe6 => s_INPUT_link_arr(0),
         probe7 => s_OUTPUT_link_arr(0)
     );
     
-----------------------------------------------------------------------------
-- Begin User_Code
-----------------------------------------------------------------------------
     
   i_Getclustertracklinker_3 : Getclustertracklinker_3
       PORT MAP (
         ap_clk => ap_clk,
         ap_rst => ap_rst,
         ap_start => ap_start,
         ap_done => ap_done,
         ap_idle => ap_idle,
         ap_ready => ap_ready,
         
         
         ClusterET_0_0_V => ClusterET_0_0_V,
         ClusterET_0_1_V => ClusterET_0_1_V,
         ClusterET_0_2_V => ClusterET_0_2_V,
         ClusterET_0_3_V => ClusterET_0_3_V,
         ClusterET_1_0_V => ClusterET_1_0_V,
         ClusterET_1_1_V => ClusterET_1_1_V,
         ClusterET_1_2_V => ClusterET_1_2_V,
         ClusterET_1_3_V => ClusterET_1_3_V,
         ClusterET_2_0_V => ClusterET_2_0_V,
         ClusterET_2_1_V => ClusterET_2_1_V,
         ClusterET_2_2_V => ClusterET_2_2_V,
         ClusterET_2_3_V => ClusterET_2_3_V,
         ClusterET_3_0_V => ClusterET_3_0_V,
         ClusterET_3_1_V => ClusterET_3_1_V,
         ClusterET_3_2_V => ClusterET_3_2_V,
         ClusterET_3_3_V => ClusterET_3_3_V,
         ClusterET_4_0_V => ClusterET_4_0_V,
         ClusterET_4_1_V => ClusterET_4_1_V,
         ClusterET_4_2_V => ClusterET_4_2_V,
         ClusterET_4_3_V => ClusterET_4_3_V,
         ClusterET_5_0_V => ClusterET_5_0_V,
         ClusterET_5_1_V => ClusterET_5_1_V,
         ClusterET_5_2_V => ClusterET_5_2_V,
         ClusterET_5_3_V => ClusterET_5_3_V,
         ClusterET_6_0_V => ClusterET_6_0_V,
         ClusterET_6_1_V => ClusterET_6_1_V,
         ClusterET_6_2_V => ClusterET_6_2_V,
         ClusterET_6_3_V => ClusterET_6_3_V,
         ClusterET_7_0_V => ClusterET_7_0_V,
         ClusterET_7_1_V => ClusterET_7_1_V,
         ClusterET_7_2_V => ClusterET_7_2_V,
         ClusterET_7_3_V => ClusterET_7_3_V,
         ClusterET_8_0_V => ClusterET_8_0_V,
         ClusterET_8_1_V => ClusterET_8_1_V,
         ClusterET_8_2_V => ClusterET_8_2_V,
         ClusterET_8_3_V => ClusterET_8_3_V,
         ClusterET_9_0_V => ClusterET_9_0_V,
         ClusterET_9_1_V => ClusterET_9_1_V,
         ClusterET_9_2_V => ClusterET_9_2_V,
         ClusterET_9_3_V => ClusterET_9_3_V,
         ClusterET_10_0_V => ClusterET_10_0_V,
         ClusterET_10_1_V => ClusterET_10_1_V,
         ClusterET_10_2_V => ClusterET_10_2_V,
         ClusterET_10_3_V => ClusterET_10_3_V,
         ClusterET_11_0_V => ClusterET_11_0_V,
         ClusterET_11_1_V => ClusterET_11_1_V,
         ClusterET_11_2_V => ClusterET_11_2_V,
         ClusterET_11_3_V => ClusterET_11_3_V,
         ClusterET_12_0_V => ClusterET_12_0_V,
         ClusterET_12_1_V => ClusterET_12_1_V,
         ClusterET_12_2_V => ClusterET_12_2_V,
         ClusterET_12_3_V => ClusterET_12_3_V,
         ClusterET_13_0_V => ClusterET_13_0_V,
         ClusterET_13_1_V => ClusterET_13_1_V,
         ClusterET_13_2_V => ClusterET_13_2_V,
         ClusterET_13_3_V => ClusterET_13_3_V,
         ClusterET_14_0_V => ClusterET_14_0_V,
         ClusterET_14_1_V => ClusterET_14_1_V,
         ClusterET_14_2_V => ClusterET_14_2_V,
         ClusterET_14_3_V => ClusterET_14_3_V,
         ClusterET_15_0_V => ClusterET_15_0_V,
         ClusterET_15_1_V => ClusterET_15_1_V,
         ClusterET_15_2_V => ClusterET_15_2_V,
         ClusterET_15_3_V => ClusterET_15_3_V,
         ClusterET_16_0_V => ClusterET_16_0_V,
         ClusterET_16_1_V => ClusterET_16_1_V,
         ClusterET_16_2_V => ClusterET_16_2_V,
         ClusterET_16_3_V => ClusterET_16_3_V,
         
         
         peakEta_0_0_V => peakEta_0_0_V,
         peakEta_0_1_V => peakEta_0_1_V,
         peakEta_0_2_V => peakEta_0_2_V,
         peakEta_0_3_V => peakEta_0_3_V,
         peakEta_1_0_V => peakEta_1_0_V,
         peakEta_1_1_V => peakEta_1_1_V,
         peakEta_1_2_V => peakEta_1_2_V,
         peakEta_1_3_V => peakEta_1_3_V,
         peakEta_2_0_V => peakEta_2_0_V,
         peakEta_2_1_V => peakEta_2_1_V,
         peakEta_2_2_V => peakEta_2_2_V,
         peakEta_2_3_V => peakEta_2_3_V,
         peakEta_3_0_V => peakEta_3_0_V,
         peakEta_3_1_V => peakEta_3_1_V,
         peakEta_3_2_V => peakEta_3_2_V,
         peakEta_3_3_V => peakEta_3_3_V,
         peakEta_4_0_V => peakEta_4_0_V,
         peakEta_4_1_V => peakEta_4_1_V,
         peakEta_4_2_V => peakEta_4_2_V,
         peakEta_4_3_V => peakEta_4_3_V,
         peakEta_5_0_V => peakEta_5_0_V,
         peakEta_5_1_V => peakEta_5_1_V,
         peakEta_5_2_V => peakEta_5_2_V,
         peakEta_5_3_V => peakEta_5_3_V,
         peakEta_6_0_V => peakEta_6_0_V,
         peakEta_6_1_V => peakEta_6_1_V,
         peakEta_6_2_V => peakEta_6_2_V,
         peakEta_6_3_V => peakEta_6_3_V,
         peakEta_7_0_V => peakEta_7_0_V,
         peakEta_7_1_V => peakEta_7_1_V,
         peakEta_7_2_V => peakEta_7_2_V,
         peakEta_7_3_V => peakEta_7_3_V,
         peakEta_8_0_V => peakEta_8_0_V,
         peakEta_8_1_V => peakEta_8_1_V,
         peakEta_8_2_V => peakEta_8_2_V,
         peakEta_8_3_V => peakEta_8_3_V,
         peakEta_9_0_V => peakEta_9_0_V,
         peakEta_9_1_V => peakEta_9_1_V,
         peakEta_9_2_V => peakEta_9_2_V,
         peakEta_9_3_V => peakEta_9_3_V,
         peakEta_10_0_V => peakEta_10_0_V,
         peakEta_10_1_V => peakEta_10_1_V,
         peakEta_10_2_V => peakEta_10_2_V,
         peakEta_10_3_V => peakEta_10_3_V,
         peakEta_11_0_V => peakEta_11_0_V,
         peakEta_11_1_V => peakEta_11_1_V,
         peakEta_11_2_V => peakEta_11_2_V,
         peakEta_11_3_V => peakEta_11_3_V,
         peakEta_12_0_V => peakEta_12_0_V,
         peakEta_12_1_V => peakEta_12_1_V,
         peakEta_12_2_V => peakEta_12_2_V,
         peakEta_12_3_V => peakEta_12_3_V,
         peakEta_13_0_V => peakEta_13_0_V,
         peakEta_13_1_V => peakEta_13_1_V,
         peakEta_13_2_V => peakEta_13_2_V,
         peakEta_13_3_V => peakEta_13_3_V,
         peakEta_14_0_V => peakEta_14_0_V,
         peakEta_14_1_V => peakEta_14_1_V,
         peakEta_14_2_V => peakEta_14_2_V,
         peakEta_14_3_V => peakEta_14_3_V,
         peakEta_15_0_V => peakEta_15_0_V,
         peakEta_15_1_V => peakEta_15_1_V,
         peakEta_15_2_V => peakEta_15_2_V,
         peakEta_15_3_V => peakEta_15_3_V,
         peakEta_16_0_V => peakEta_16_0_V,
         peakEta_16_1_V => peakEta_16_1_V,
         peakEta_16_2_V => peakEta_16_2_V,
         peakEta_16_3_V => peakEta_16_3_V,
         
         
         peakPhi_0_0_V => peakPhi_0_0_V,
         peakPhi_0_1_V => peakPhi_0_1_V,
         peakPhi_0_2_V => peakPhi_0_2_V,
         peakPhi_0_3_V => peakPhi_0_3_V,
         peakPhi_1_0_V => peakPhi_1_0_V,
         peakPhi_1_1_V => peakPhi_1_1_V,
         peakPhi_1_2_V => peakPhi_1_2_V,
         peakPhi_1_3_V => peakPhi_1_3_V,
         peakPhi_2_0_V => peakPhi_2_0_V,
         peakPhi_2_1_V => peakPhi_2_1_V,
         peakPhi_2_2_V => peakPhi_2_2_V,
         peakPhi_2_3_V => peakPhi_2_3_V,
         peakPhi_3_0_V => peakPhi_3_0_V,
         peakPhi_3_1_V => peakPhi_3_1_V,
         peakPhi_3_2_V => peakPhi_3_2_V,
         peakPhi_3_3_V => peakPhi_3_3_V,
         peakPhi_4_0_V => peakPhi_4_0_V,
         peakPhi_4_1_V => peakPhi_4_1_V,
         peakPhi_4_2_V => peakPhi_4_2_V,
         peakPhi_4_3_V => peakPhi_4_3_V,
         peakPhi_5_0_V => peakPhi_5_0_V,
         peakPhi_5_1_V => peakPhi_5_1_V,
         peakPhi_5_2_V => peakPhi_5_2_V,
         peakPhi_5_3_V => peakPhi_5_3_V,
         peakPhi_6_0_V => peakPhi_6_0_V,
         peakPhi_6_1_V => peakPhi_6_1_V,
         peakPhi_6_2_V => peakPhi_6_2_V,
         peakPhi_6_3_V => peakPhi_6_3_V,
         peakPhi_7_0_V => peakPhi_7_0_V,
         peakPhi_7_1_V => peakPhi_7_1_V,
         peakPhi_7_2_V => peakPhi_7_2_V,
         peakPhi_7_3_V => peakPhi_7_3_V,
         peakPhi_8_0_V => peakPhi_8_0_V,
         peakPhi_8_1_V => peakPhi_8_1_V,
         peakPhi_8_2_V => peakPhi_8_2_V,
         peakPhi_8_3_V => peakPhi_8_3_V,
         peakPhi_9_0_V => peakPhi_9_0_V,
         peakPhi_9_1_V => peakPhi_9_1_V,
         peakPhi_9_2_V => peakPhi_9_2_V,
         peakPhi_9_3_V => peakPhi_9_3_V,
         peakPhi_10_0_V => peakPhi_10_0_V,
         peakPhi_10_1_V => peakPhi_10_1_V,
         peakPhi_10_2_V => peakPhi_10_2_V,
         peakPhi_10_3_V => peakPhi_10_3_V,
         peakPhi_11_0_V => peakPhi_11_0_V,
         peakPhi_11_1_V => peakPhi_11_1_V,
         peakPhi_11_2_V => peakPhi_11_2_V,
         peakPhi_11_3_V => peakPhi_11_3_V,
         peakPhi_12_0_V => peakPhi_12_0_V,
         peakPhi_12_1_V => peakPhi_12_1_V,
         peakPhi_12_2_V => peakPhi_12_2_V,
         peakPhi_12_3_V => peakPhi_12_3_V,
         peakPhi_13_0_V => peakPhi_13_0_V,
         peakPhi_13_1_V => peakPhi_13_1_V,
         peakPhi_13_2_V => peakPhi_13_2_V,
         peakPhi_13_3_V => peakPhi_13_3_V,
         peakPhi_14_0_V => peakPhi_14_0_V,
         peakPhi_14_1_V => peakPhi_14_1_V,
         peakPhi_14_2_V => peakPhi_14_2_V,
         peakPhi_14_3_V => peakPhi_14_3_V,
         peakPhi_15_0_V => peakPhi_15_0_V,
         peakPhi_15_1_V => peakPhi_15_1_V,
         peakPhi_15_2_V => peakPhi_15_2_V,
         peakPhi_15_3_V => peakPhi_15_3_V,
         peakPhi_16_0_V => peakPhi_16_0_V,
         peakPhi_16_1_V => peakPhi_16_1_V,
         peakPhi_16_2_V => peakPhi_16_2_V,
         peakPhi_16_3_V => peakPhi_16_3_V,
         
         
         trackPT_0_V => trackPT_0_V,
         trackPT_1_V => trackPT_1_V,
         trackPT_2_V => trackPT_2_V,
         trackPT_3_V => trackPT_3_V,
         trackPT_4_V => trackPT_4_V,
         trackPT_5_V => trackPT_5_V,
         trackPT_6_V => trackPT_6_V,
         trackPT_7_V => trackPT_7_V,
         trackPT_8_V => trackPT_8_V,
         trackPT_9_V => trackPT_9_V,
         
         
         trackEta_0_V => trackEta_0_V,
         trackEta_1_V => trackEta_1_V,
         trackEta_2_V => trackEta_2_V,
         trackEta_3_V => trackEta_3_V,
         trackEta_4_V => trackEta_4_V,
         trackEta_5_V => trackEta_5_V,
         trackEta_6_V => trackEta_6_V,
         trackEta_7_V => trackEta_7_V,
         trackEta_8_V => trackEta_8_V,
         trackEta_9_V => trackEta_9_V,
         
         
         trackPhi_0_V => trackPhi_0_V,
         trackPhi_1_V => trackPhi_1_V,
         trackPhi_2_V => trackPhi_2_V,
         trackPhi_3_V => trackPhi_3_V,
         trackPhi_4_V => trackPhi_4_V,
         trackPhi_5_V => trackPhi_5_V,
         trackPhi_6_V => trackPhi_6_V,
         trackPhi_7_V => trackPhi_7_V,
         trackPhi_8_V => trackPhi_8_V,
         trackPhi_9_V => trackPhi_9_V,
         
         
         output_linkedTrackPT_0_V => output_linkedTrackPT_0_V,
         output_linkedTrackPT_1_V => output_linkedTrackPT_1_V,
         output_linkedTrackPT_2_V => output_linkedTrackPT_2_V,
         output_linkedTrackPT_3_V => output_linkedTrackPT_3_V,
         output_linkedTrackPT_4_V => output_linkedTrackPT_4_V,
         output_linkedTrackPT_5_V => output_linkedTrackPT_5_V,
         output_linkedTrackPT_6_V => output_linkedTrackPT_6_V,
         output_linkedTrackPT_7_V => output_linkedTrackPT_7_V,
         output_linkedTrackPT_8_V => output_linkedTrackPT_8_V,
         output_linkedTrackPT_9_V => output_linkedTrackPT_9_V,
         
         
         output_linkedTrackEta_0_V => output_linkedTrackEta_0_V,
         output_linkedTrackEta_1_V => output_linkedTrackEta_1_V,
         output_linkedTrackEta_2_V => output_linkedTrackEta_2_V,
         output_linkedTrackEta_3_V => output_linkedTrackEta_3_V,
         output_linkedTrackEta_4_V => output_linkedTrackEta_4_V,
         output_linkedTrackEta_5_V => output_linkedTrackEta_5_V,
         output_linkedTrackEta_6_V => output_linkedTrackEta_6_V,
         output_linkedTrackEta_7_V => output_linkedTrackEta_7_V,
         output_linkedTrackEta_8_V => output_linkedTrackEta_8_V,
         output_linkedTrackEta_9_V => output_linkedTrackEta_9_V,
         
         
         output_linkedTrackPhi_0_V => output_linkedTrackPhi_0_V,
         output_linkedTrackPhi_1_V => output_linkedTrackPhi_1_V,
         output_linkedTrackPhi_2_V => output_linkedTrackPhi_2_V,
         output_linkedTrackPhi_3_V => output_linkedTrackPhi_3_V,
         output_linkedTrackPhi_4_V => output_linkedTrackPhi_4_V,
         output_linkedTrackPhi_5_V => output_linkedTrackPhi_5_V,
         output_linkedTrackPhi_6_V => output_linkedTrackPhi_6_V,
         output_linkedTrackPhi_7_V => output_linkedTrackPhi_7_V,
         output_linkedTrackPhi_8_V => output_linkedTrackPhi_8_V,
         output_linkedTrackPhi_9_V => output_linkedTrackPhi_9_V,
         
         
         output_linkedTrackQuality_0_V => output_linkedTrackQuality_0_V,
         output_linkedTrackQuality_1_V => output_linkedTrackQuality_1_V,
         output_linkedTrackQuality_2_V => output_linkedTrackQuality_2_V,
         output_linkedTrackQuality_3_V => output_linkedTrackQuality_3_V,
         output_linkedTrackQuality_4_V => output_linkedTrackQuality_4_V,
         output_linkedTrackQuality_5_V => output_linkedTrackQuality_5_V,
         output_linkedTrackQuality_6_V => output_linkedTrackQuality_6_V,
         output_linkedTrackQuality_7_V => output_linkedTrackQuality_7_V,
         output_linkedTrackQuality_8_V => output_linkedTrackQuality_8_V,
         output_linkedTrackQuality_9_V => output_linkedTrackQuality_9_V,
         
         
         output_neutralClusterET_0_V => output_neutralClusterET_0_V,
         output_neutralClusterET_1_V => output_neutralClusterET_1_V,
         output_neutralClusterET_2_V => output_neutralClusterET_2_V,
         output_neutralClusterET_3_V => output_neutralClusterET_3_V,
         output_neutralClusterET_4_V => output_neutralClusterET_4_V,
         output_neutralClusterET_5_V => output_neutralClusterET_5_V,
         output_neutralClusterET_6_V => output_neutralClusterET_6_V,
         output_neutralClusterET_7_V => output_neutralClusterET_7_V,
         output_neutralClusterET_8_V => output_neutralClusterET_8_V,
         output_neutralClusterET_9_V => output_neutralClusterET_9_V,
         output_neutralClusterET_10_V => output_neutralClusterET_10_V,
         output_neutralClusterET_11_V => output_neutralClusterET_11_V,
         output_neutralClusterET_12_V => output_neutralClusterET_12_V,
         output_neutralClusterET_13_V => output_neutralClusterET_13_V,
         output_neutralClusterET_14_V => output_neutralClusterET_14_V,
         output_neutralClusterET_15_V => output_neutralClusterET_15_V,
         output_neutralClusterET_16_V => output_neutralClusterET_16_V,
         output_neutralClusterET_17_V => output_neutralClusterET_17_V,
         output_neutralClusterET_18_V => output_neutralClusterET_18_V,
         output_neutralClusterET_19_V => output_neutralClusterET_19_V,
         output_neutralClusterET_20_V => output_neutralClusterET_20_V,
         output_neutralClusterET_21_V => output_neutralClusterET_21_V,
         output_neutralClusterET_22_V => output_neutralClusterET_22_V,
         output_neutralClusterET_23_V => output_neutralClusterET_23_V,
         output_neutralClusterET_24_V => output_neutralClusterET_24_V,
         output_neutralClusterET_25_V => output_neutralClusterET_25_V,
         output_neutralClusterET_26_V => output_neutralClusterET_26_V,
         output_neutralClusterET_27_V => output_neutralClusterET_27_V,
         output_neutralClusterET_28_V => output_neutralClusterET_28_V,
         output_neutralClusterET_29_V => output_neutralClusterET_29_V,
         output_neutralClusterET_30_V => output_neutralClusterET_30_V,
         output_neutralClusterET_31_V => output_neutralClusterET_31_V,
         output_neutralClusterET_32_V => output_neutralClusterET_32_V,
         output_neutralClusterET_33_V => output_neutralClusterET_33_V,
         output_neutralClusterET_34_V => output_neutralClusterET_34_V,
         output_neutralClusterET_35_V => output_neutralClusterET_35_V,
         output_neutralClusterET_36_V => output_neutralClusterET_36_V,
         output_neutralClusterET_37_V => output_neutralClusterET_37_V,
         output_neutralClusterET_38_V => output_neutralClusterET_38_V,
         output_neutralClusterET_39_V => output_neutralClusterET_39_V,
         output_neutralClusterET_40_V => output_neutralClusterET_40_V,
         output_neutralClusterET_41_V => output_neutralClusterET_41_V,
         output_neutralClusterET_42_V => output_neutralClusterET_42_V,
         output_neutralClusterET_43_V => output_neutralClusterET_43_V,
         output_neutralClusterET_44_V => output_neutralClusterET_44_V,
         output_neutralClusterET_45_V => output_neutralClusterET_45_V,
         output_neutralClusterET_46_V => output_neutralClusterET_46_V,
         output_neutralClusterET_47_V => output_neutralClusterET_47_V,
         output_neutralClusterET_48_V => output_neutralClusterET_48_V,
         output_neutralClusterET_49_V => output_neutralClusterET_49_V,
         output_neutralClusterET_50_V => output_neutralClusterET_50_V,
         output_neutralClusterET_51_V => output_neutralClusterET_51_V,
         output_neutralClusterET_52_V => output_neutralClusterET_52_V,
         output_neutralClusterET_53_V => output_neutralClusterET_53_V,
         output_neutralClusterET_54_V => output_neutralClusterET_54_V,
         output_neutralClusterET_55_V => output_neutralClusterET_55_V,
         output_neutralClusterET_56_V => output_neutralClusterET_56_V,
         output_neutralClusterET_57_V => output_neutralClusterET_57_V,
         output_neutralClusterET_58_V => output_neutralClusterET_58_V,
         output_neutralClusterET_59_V => output_neutralClusterET_59_V,
         output_neutralClusterET_60_V => output_neutralClusterET_60_V,
         output_neutralClusterET_61_V => output_neutralClusterET_61_V,
         output_neutralClusterET_62_V => output_neutralClusterET_62_V,
         output_neutralClusterET_63_V => output_neutralClusterET_63_V,
         output_neutralClusterET_64_V => output_neutralClusterET_64_V,
         output_neutralClusterET_65_V => output_neutralClusterET_65_V,
         output_neutralClusterET_66_V => output_neutralClusterET_66_V,
         output_neutralClusterET_67_V => output_neutralClusterET_67_V,
         
         
         output_neutralClusterEta_0_V => output_neutralClusterEta_0_V,
         output_neutralClusterEta_1_V => output_neutralClusterEta_1_V,
         output_neutralClusterEta_2_V => output_neutralClusterEta_2_V,
         output_neutralClusterEta_3_V => output_neutralClusterEta_3_V,
         output_neutralClusterEta_4_V => output_neutralClusterEta_4_V,
         output_neutralClusterEta_5_V => output_neutralClusterEta_5_V,
         output_neutralClusterEta_6_V => output_neutralClusterEta_6_V,
         output_neutralClusterEta_7_V => output_neutralClusterEta_7_V,
         output_neutralClusterEta_8_V => output_neutralClusterEta_8_V,
         output_neutralClusterEta_9_V => output_neutralClusterEta_9_V,
         output_neutralClusterEta_10_V => output_neutralClusterEta_10_V,
         output_neutralClusterEta_11_V => output_neutralClusterEta_11_V,
         output_neutralClusterEta_12_V => output_neutralClusterEta_12_V,
         output_neutralClusterEta_13_V => output_neutralClusterEta_13_V,
         output_neutralClusterEta_14_V => output_neutralClusterEta_14_V,
         output_neutralClusterEta_15_V => output_neutralClusterEta_15_V,
         output_neutralClusterEta_16_V => output_neutralClusterEta_16_V,
         output_neutralClusterEta_17_V => output_neutralClusterEta_17_V,
         output_neutralClusterEta_18_V => output_neutralClusterEta_18_V,
         output_neutralClusterEta_19_V => output_neutralClusterEta_19_V,
         output_neutralClusterEta_20_V => output_neutralClusterEta_20_V,
         output_neutralClusterEta_21_V => output_neutralClusterEta_21_V,
         output_neutralClusterEta_22_V => output_neutralClusterEta_22_V,
         output_neutralClusterEta_23_V => output_neutralClusterEta_23_V,
         output_neutralClusterEta_24_V => output_neutralClusterEta_24_V,
         output_neutralClusterEta_25_V => output_neutralClusterEta_25_V,
         output_neutralClusterEta_26_V => output_neutralClusterEta_26_V,
         output_neutralClusterEta_27_V => output_neutralClusterEta_27_V,
         output_neutralClusterEta_28_V => output_neutralClusterEta_28_V,
         output_neutralClusterEta_29_V => output_neutralClusterEta_29_V,
         output_neutralClusterEta_30_V => output_neutralClusterEta_30_V,
         output_neutralClusterEta_31_V => output_neutralClusterEta_31_V,
         output_neutralClusterEta_32_V => output_neutralClusterEta_32_V,
         output_neutralClusterEta_33_V => output_neutralClusterEta_33_V,
         output_neutralClusterEta_34_V => output_neutralClusterEta_34_V,
         output_neutralClusterEta_35_V => output_neutralClusterEta_35_V,
         output_neutralClusterEta_36_V => output_neutralClusterEta_36_V,
         output_neutralClusterEta_37_V => output_neutralClusterEta_37_V,
         output_neutralClusterEta_38_V => output_neutralClusterEta_38_V,
         output_neutralClusterEta_39_V => output_neutralClusterEta_39_V,
         output_neutralClusterEta_40_V => output_neutralClusterEta_40_V,
         output_neutralClusterEta_41_V => output_neutralClusterEta_41_V,
         output_neutralClusterEta_42_V => output_neutralClusterEta_42_V,
         output_neutralClusterEta_43_V => output_neutralClusterEta_43_V,
         output_neutralClusterEta_44_V => output_neutralClusterEta_44_V,
         output_neutralClusterEta_45_V => output_neutralClusterEta_45_V,
         output_neutralClusterEta_46_V => output_neutralClusterEta_46_V,
         output_neutralClusterEta_47_V => output_neutralClusterEta_47_V,
         output_neutralClusterEta_48_V => output_neutralClusterEta_48_V,
         output_neutralClusterEta_49_V => output_neutralClusterEta_49_V,
         output_neutralClusterEta_50_V => output_neutralClusterEta_50_V,
         output_neutralClusterEta_51_V => output_neutralClusterEta_51_V,
         output_neutralClusterEta_52_V => output_neutralClusterEta_52_V,
         output_neutralClusterEta_53_V => output_neutralClusterEta_53_V,
         output_neutralClusterEta_54_V => output_neutralClusterEta_54_V,
         output_neutralClusterEta_55_V => output_neutralClusterEta_55_V,
         output_neutralClusterEta_56_V => output_neutralClusterEta_56_V,
         output_neutralClusterEta_57_V => output_neutralClusterEta_57_V,
         output_neutralClusterEta_58_V => output_neutralClusterEta_58_V,
         output_neutralClusterEta_59_V => output_neutralClusterEta_59_V,
         output_neutralClusterEta_60_V => output_neutralClusterEta_60_V,
         output_neutralClusterEta_61_V => output_neutralClusterEta_61_V,
         output_neutralClusterEta_62_V => output_neutralClusterEta_62_V,
         output_neutralClusterEta_63_V => output_neutralClusterEta_63_V,
         output_neutralClusterEta_64_V => output_neutralClusterEta_64_V,
         output_neutralClusterEta_65_V => output_neutralClusterEta_65_V,
         output_neutralClusterEta_66_V => output_neutralClusterEta_66_V,
         output_neutralClusterEta_67_V => output_neutralClusterEta_67_V,
         
         
         output_neutralClusterPhi_0_V => output_neutralClusterPhi_0_V,
         output_neutralClusterPhi_1_V => output_neutralClusterPhi_1_V,
         output_neutralClusterPhi_2_V => output_neutralClusterPhi_2_V,
         output_neutralClusterPhi_3_V => output_neutralClusterPhi_3_V,
         output_neutralClusterPhi_4_V => output_neutralClusterPhi_4_V,
         output_neutralClusterPhi_5_V => output_neutralClusterPhi_5_V,
         output_neutralClusterPhi_6_V => output_neutralClusterPhi_6_V,
         output_neutralClusterPhi_7_V => output_neutralClusterPhi_7_V,
         output_neutralClusterPhi_8_V => output_neutralClusterPhi_8_V,
         output_neutralClusterPhi_9_V => output_neutralClusterPhi_9_V,
         output_neutralClusterPhi_10_V => output_neutralClusterPhi_10_V,
         output_neutralClusterPhi_11_V => output_neutralClusterPhi_11_V,
         output_neutralClusterPhi_12_V => output_neutralClusterPhi_12_V,
         output_neutralClusterPhi_13_V => output_neutralClusterPhi_13_V,
         output_neutralClusterPhi_14_V => output_neutralClusterPhi_14_V,
         output_neutralClusterPhi_15_V => output_neutralClusterPhi_15_V,
         output_neutralClusterPhi_16_V => output_neutralClusterPhi_16_V,
         output_neutralClusterPhi_17_V => output_neutralClusterPhi_17_V,
         output_neutralClusterPhi_18_V => output_neutralClusterPhi_18_V,
         output_neutralClusterPhi_19_V => output_neutralClusterPhi_19_V,
         output_neutralClusterPhi_20_V => output_neutralClusterPhi_20_V,
         output_neutralClusterPhi_21_V => output_neutralClusterPhi_21_V,
         output_neutralClusterPhi_22_V => output_neutralClusterPhi_22_V,
         output_neutralClusterPhi_23_V => output_neutralClusterPhi_23_V,
         output_neutralClusterPhi_24_V => output_neutralClusterPhi_24_V,
         output_neutralClusterPhi_25_V => output_neutralClusterPhi_25_V,
         output_neutralClusterPhi_26_V => output_neutralClusterPhi_26_V,
         output_neutralClusterPhi_27_V => output_neutralClusterPhi_27_V,
         output_neutralClusterPhi_28_V => output_neutralClusterPhi_28_V,
         output_neutralClusterPhi_29_V => output_neutralClusterPhi_29_V,
         output_neutralClusterPhi_30_V => output_neutralClusterPhi_30_V,
         output_neutralClusterPhi_31_V => output_neutralClusterPhi_31_V,
         output_neutralClusterPhi_32_V => output_neutralClusterPhi_32_V,
         output_neutralClusterPhi_33_V => output_neutralClusterPhi_33_V,
         output_neutralClusterPhi_34_V => output_neutralClusterPhi_34_V,
         output_neutralClusterPhi_35_V => output_neutralClusterPhi_35_V,
         output_neutralClusterPhi_36_V => output_neutralClusterPhi_36_V,
         output_neutralClusterPhi_37_V => output_neutralClusterPhi_37_V,
         output_neutralClusterPhi_38_V => output_neutralClusterPhi_38_V,
         output_neutralClusterPhi_39_V => output_neutralClusterPhi_39_V,
         output_neutralClusterPhi_40_V => output_neutralClusterPhi_40_V,
         output_neutralClusterPhi_41_V => output_neutralClusterPhi_41_V,
         output_neutralClusterPhi_42_V => output_neutralClusterPhi_42_V,
         output_neutralClusterPhi_43_V => output_neutralClusterPhi_43_V,
         output_neutralClusterPhi_44_V => output_neutralClusterPhi_44_V,
         output_neutralClusterPhi_45_V => output_neutralClusterPhi_45_V,
         output_neutralClusterPhi_46_V => output_neutralClusterPhi_46_V,
         output_neutralClusterPhi_47_V => output_neutralClusterPhi_47_V,
         output_neutralClusterPhi_48_V => output_neutralClusterPhi_48_V,
         output_neutralClusterPhi_49_V => output_neutralClusterPhi_49_V,
         output_neutralClusterPhi_50_V => output_neutralClusterPhi_50_V,
         output_neutralClusterPhi_51_V => output_neutralClusterPhi_51_V,
         output_neutralClusterPhi_52_V => output_neutralClusterPhi_52_V,
         output_neutralClusterPhi_53_V => output_neutralClusterPhi_53_V,
         output_neutralClusterPhi_54_V => output_neutralClusterPhi_54_V,
         output_neutralClusterPhi_55_V => output_neutralClusterPhi_55_V,
         output_neutralClusterPhi_56_V => output_neutralClusterPhi_56_V,
         output_neutralClusterPhi_57_V => output_neutralClusterPhi_57_V,
         output_neutralClusterPhi_58_V => output_neutralClusterPhi_58_V,
         output_neutralClusterPhi_59_V => output_neutralClusterPhi_59_V,
         output_neutralClusterPhi_60_V => output_neutralClusterPhi_60_V,
         output_neutralClusterPhi_61_V => output_neutralClusterPhi_61_V,
         output_neutralClusterPhi_62_V => output_neutralClusterPhi_62_V,
         output_neutralClusterPhi_63_V => output_neutralClusterPhi_63_V,
         output_neutralClusterPhi_64_V => output_neutralClusterPhi_64_V,
         output_neutralClusterPhi_65_V => output_neutralClusterPhi_65_V,
         output_neutralClusterPhi_66_V => output_neutralClusterPhi_66_V,
         output_neutralClusterPhi_67_V => output_neutralClusterPhi_67_V
         
       );

-----------------------------------------------------------------------------
-- Configuration registers              
   
-----------------------------------------------------------------------------

-- Input and Output Links

ClusterET_0_0_V <= s_INPUT_LINK_ARR( 0 )(9 downto 0);
peakEta_0_0_V <= s_INPUT_LINK_ARR( 0 )(12 downto 10);
peakPhi_0_0_V <= s_INPUT_LINK_ARR( 0 )(15 downto 13);
ClusterET_0_1_V <= s_INPUT_LINK_ARR( 0 )(25 downto 16);
peakEta_0_1_V <= s_INPUT_LINK_ARR( 0 )(28 downto 26);
peakPhi_0_1_V <= s_INPUT_LINK_ARR( 0 )(31 downto 29);
ClusterET_0_2_V <= s_INPUT_LINK_ARR( 0 )(41 downto 32);
peakEta_0_2_V <= s_INPUT_LINK_ARR( 0 )(44 downto 42);
peakPhi_0_2_V <= s_INPUT_LINK_ARR( 0 )(47 downto 45);
ClusterET_0_3_V <= s_INPUT_LINK_ARR( 0 )(57 downto 48);
peakEta_0_3_V <= s_INPUT_LINK_ARR( 0 )(60 downto 58);
peakPhi_0_3_V <= s_INPUT_LINK_ARR( 0 )(63 downto 61);
ClusterET_1_0_V <= s_INPUT_LINK_ARR( 0 )(73 downto 64);
peakEta_1_0_V <= s_INPUT_LINK_ARR( 0 )(76 downto 74);
peakPhi_1_0_V <= s_INPUT_LINK_ARR( 0 )(79 downto 77);
ClusterET_1_1_V <= s_INPUT_LINK_ARR( 0 )(89 downto 80);
peakEta_1_1_V <= s_INPUT_LINK_ARR( 0 )(92 downto 90);
peakPhi_1_1_V <= s_INPUT_LINK_ARR( 0 )(95 downto 93);
ClusterET_1_2_V <= s_INPUT_LINK_ARR( 0 )(105 downto 96);
peakEta_1_2_V <= s_INPUT_LINK_ARR( 0 )(108 downto 106);
peakPhi_1_2_V <= s_INPUT_LINK_ARR( 0 )(111 downto 109);
ClusterET_1_3_V <= s_INPUT_LINK_ARR( 0 )(121 downto 112);
peakEta_1_3_V <= s_INPUT_LINK_ARR( 0 )(124 downto 122);
peakPhi_1_3_V <= s_INPUT_LINK_ARR( 0 )(127 downto 125);
ClusterET_2_0_V <= s_INPUT_LINK_ARR( 0 )(137 downto 128);
peakEta_2_0_V <= s_INPUT_LINK_ARR( 0 )(140 downto 138);
peakPhi_2_0_V <= s_INPUT_LINK_ARR( 0 )(143 downto 141);
ClusterET_2_1_V <= s_INPUT_LINK_ARR( 0 )(153 downto 144);
peakEta_2_1_V <= s_INPUT_LINK_ARR( 0 )(156 downto 154);
peakPhi_2_1_V <= s_INPUT_LINK_ARR( 0 )(159 downto 157);
ClusterET_2_2_V <= s_INPUT_LINK_ARR( 0 )(169 downto 160);
peakEta_2_2_V <= s_INPUT_LINK_ARR( 0 )(172 downto 170);
peakPhi_2_2_V <= s_INPUT_LINK_ARR( 0 )(175 downto 173);
ClusterET_2_3_V <= s_INPUT_LINK_ARR( 0 )(185 downto 176);
peakEta_2_3_V <= s_INPUT_LINK_ARR( 0 )(188 downto 186);
peakPhi_2_3_V <= s_INPUT_LINK_ARR( 0 )(191 downto 189);
ClusterET_3_0_V <= s_INPUT_LINK_ARR( 1 )(9 downto 0);
peakEta_3_0_V <= s_INPUT_LINK_ARR( 1 )(12 downto 10);
peakPhi_3_0_V <= s_INPUT_LINK_ARR( 1 )(15 downto 13);
ClusterET_3_1_V <= s_INPUT_LINK_ARR( 1 )(25 downto 16);
peakEta_3_1_V <= s_INPUT_LINK_ARR( 1 )(28 downto 26);
peakPhi_3_1_V <= s_INPUT_LINK_ARR( 1 )(31 downto 29);
ClusterET_3_2_V <= s_INPUT_LINK_ARR( 1 )(41 downto 32);
peakEta_3_2_V <= s_INPUT_LINK_ARR( 1 )(44 downto 42);
peakPhi_3_2_V <= s_INPUT_LINK_ARR( 1 )(47 downto 45);
ClusterET_3_3_V <= s_INPUT_LINK_ARR( 1 )(57 downto 48);
peakEta_3_3_V <= s_INPUT_LINK_ARR( 1 )(60 downto 58);
peakPhi_3_3_V <= s_INPUT_LINK_ARR( 1 )(63 downto 61);
ClusterET_4_0_V <= s_INPUT_LINK_ARR( 1 )(73 downto 64);
peakEta_4_0_V <= s_INPUT_LINK_ARR( 1 )(76 downto 74);
peakPhi_4_0_V <= s_INPUT_LINK_ARR( 1 )(79 downto 77);
ClusterET_4_1_V <= s_INPUT_LINK_ARR( 1 )(89 downto 80);
peakEta_4_1_V <= s_INPUT_LINK_ARR( 1 )(92 downto 90);
peakPhi_4_1_V <= s_INPUT_LINK_ARR( 1 )(95 downto 93);
ClusterET_4_2_V <= s_INPUT_LINK_ARR( 1 )(105 downto 96);
peakEta_4_2_V <= s_INPUT_LINK_ARR( 1 )(108 downto 106);
peakPhi_4_2_V <= s_INPUT_LINK_ARR( 1 )(111 downto 109);
ClusterET_4_3_V <= s_INPUT_LINK_ARR( 1 )(121 downto 112);
peakEta_4_3_V <= s_INPUT_LINK_ARR( 1 )(124 downto 122);
peakPhi_4_3_V <= s_INPUT_LINK_ARR( 1 )(127 downto 125);
ClusterET_5_0_V <= s_INPUT_LINK_ARR( 1 )(137 downto 128);
peakEta_5_0_V <= s_INPUT_LINK_ARR( 1 )(140 downto 138);
peakPhi_5_0_V <= s_INPUT_LINK_ARR( 1 )(143 downto 141);
ClusterET_5_1_V <= s_INPUT_LINK_ARR( 1 )(153 downto 144);
peakEta_5_1_V <= s_INPUT_LINK_ARR( 1 )(156 downto 154);
peakPhi_5_1_V <= s_INPUT_LINK_ARR( 1 )(159 downto 157);
ClusterET_5_2_V <= s_INPUT_LINK_ARR( 1 )(169 downto 160);
peakEta_5_2_V <= s_INPUT_LINK_ARR( 1 )(172 downto 170);
peakPhi_5_2_V <= s_INPUT_LINK_ARR( 1 )(175 downto 173);
ClusterET_5_3_V <= s_INPUT_LINK_ARR( 1 )(185 downto 176);
peakEta_5_3_V <= s_INPUT_LINK_ARR( 1 )(188 downto 186);
peakPhi_5_3_V <= s_INPUT_LINK_ARR( 1 )(191 downto 189);
ClusterET_6_0_V <= s_INPUT_LINK_ARR( 2 )(9 downto 0);
peakEta_6_0_V <= s_INPUT_LINK_ARR( 2 )(12 downto 10);
peakPhi_6_0_V <= s_INPUT_LINK_ARR( 2 )(15 downto 13);
ClusterET_6_1_V <= s_INPUT_LINK_ARR( 2 )(25 downto 16);
peakEta_6_1_V <= s_INPUT_LINK_ARR( 2 )(28 downto 26);
peakPhi_6_1_V <= s_INPUT_LINK_ARR( 2 )(31 downto 29);
ClusterET_6_2_V <= s_INPUT_LINK_ARR( 2 )(41 downto 32);
peakEta_6_2_V <= s_INPUT_LINK_ARR( 2 )(44 downto 42);
peakPhi_6_2_V <= s_INPUT_LINK_ARR( 2 )(47 downto 45);
ClusterET_6_3_V <= s_INPUT_LINK_ARR( 2 )(57 downto 48);
peakEta_6_3_V <= s_INPUT_LINK_ARR( 2 )(60 downto 58);
peakPhi_6_3_V <= s_INPUT_LINK_ARR( 2 )(63 downto 61);
ClusterET_7_0_V <= s_INPUT_LINK_ARR( 2 )(73 downto 64);
peakEta_7_0_V <= s_INPUT_LINK_ARR( 2 )(76 downto 74);
peakPhi_7_0_V <= s_INPUT_LINK_ARR( 2 )(79 downto 77);
ClusterET_7_1_V <= s_INPUT_LINK_ARR( 2 )(89 downto 80);
peakEta_7_1_V <= s_INPUT_LINK_ARR( 2 )(92 downto 90);
peakPhi_7_1_V <= s_INPUT_LINK_ARR( 2 )(95 downto 93);
ClusterET_7_2_V <= s_INPUT_LINK_ARR( 2 )(105 downto 96);
peakEta_7_2_V <= s_INPUT_LINK_ARR( 2 )(108 downto 106);
peakPhi_7_2_V <= s_INPUT_LINK_ARR( 2 )(111 downto 109);
ClusterET_7_3_V <= s_INPUT_LINK_ARR( 2 )(121 downto 112);
peakEta_7_3_V <= s_INPUT_LINK_ARR( 2 )(124 downto 122);
peakPhi_7_3_V <= s_INPUT_LINK_ARR( 2 )(127 downto 125);
ClusterET_8_0_V <= s_INPUT_LINK_ARR( 2 )(137 downto 128);
peakEta_8_0_V <= s_INPUT_LINK_ARR( 2 )(140 downto 138);
peakPhi_8_0_V <= s_INPUT_LINK_ARR( 2 )(143 downto 141);
ClusterET_8_1_V <= s_INPUT_LINK_ARR( 2 )(153 downto 144);
peakEta_8_1_V <= s_INPUT_LINK_ARR( 2 )(156 downto 154);
peakPhi_8_1_V <= s_INPUT_LINK_ARR( 2 )(159 downto 157);
ClusterET_8_2_V <= s_INPUT_LINK_ARR( 2 )(169 downto 160);
peakEta_8_2_V <= s_INPUT_LINK_ARR( 2 )(172 downto 170);
peakPhi_8_2_V <= s_INPUT_LINK_ARR( 2 )(175 downto 173);
ClusterET_8_3_V <= s_INPUT_LINK_ARR( 2 )(185 downto 176);
peakEta_8_3_V <= s_INPUT_LINK_ARR( 2 )(188 downto 186);
peakPhi_8_3_V <= s_INPUT_LINK_ARR( 2 )(191 downto 189);
ClusterET_9_0_V <= s_INPUT_LINK_ARR( 3 )(9 downto 0);
peakEta_9_0_V <= s_INPUT_LINK_ARR( 3 )(12 downto 10);
peakPhi_9_0_V <= s_INPUT_LINK_ARR( 3 )(15 downto 13);
ClusterET_9_1_V <= s_INPUT_LINK_ARR( 3 )(25 downto 16);
peakEta_9_1_V <= s_INPUT_LINK_ARR( 3 )(28 downto 26);
peakPhi_9_1_V <= s_INPUT_LINK_ARR( 3 )(31 downto 29);
ClusterET_9_2_V <= s_INPUT_LINK_ARR( 3 )(41 downto 32);
peakEta_9_2_V <= s_INPUT_LINK_ARR( 3 )(44 downto 42);
peakPhi_9_2_V <= s_INPUT_LINK_ARR( 3 )(47 downto 45);
ClusterET_9_3_V <= s_INPUT_LINK_ARR( 3 )(57 downto 48);
peakEta_9_3_V <= s_INPUT_LINK_ARR( 3 )(60 downto 58);
peakPhi_9_3_V <= s_INPUT_LINK_ARR( 3 )(63 downto 61);
ClusterET_10_0_V <= s_INPUT_LINK_ARR( 3 )(73 downto 64);
peakEta_10_0_V <= s_INPUT_LINK_ARR( 3 )(76 downto 74);
peakPhi_10_0_V <= s_INPUT_LINK_ARR( 3 )(79 downto 77);
ClusterET_10_1_V <= s_INPUT_LINK_ARR( 3 )(89 downto 80);
peakEta_10_1_V <= s_INPUT_LINK_ARR( 3 )(92 downto 90);
peakPhi_10_1_V <= s_INPUT_LINK_ARR( 3 )(95 downto 93);
ClusterET_10_2_V <= s_INPUT_LINK_ARR( 3 )(105 downto 96);
peakEta_10_2_V <= s_INPUT_LINK_ARR( 3 )(108 downto 106);
peakPhi_10_2_V <= s_INPUT_LINK_ARR( 3 )(111 downto 109);
ClusterET_10_3_V <= s_INPUT_LINK_ARR( 3 )(121 downto 112);
peakEta_10_3_V <= s_INPUT_LINK_ARR( 3 )(124 downto 122);
peakPhi_10_3_V <= s_INPUT_LINK_ARR( 3 )(127 downto 125);
ClusterET_11_0_V <= s_INPUT_LINK_ARR( 3 )(137 downto 128);
peakEta_11_0_V <= s_INPUT_LINK_ARR( 3 )(140 downto 138);
peakPhi_11_0_V <= s_INPUT_LINK_ARR( 3 )(143 downto 141);
ClusterET_11_1_V <= s_INPUT_LINK_ARR( 3 )(153 downto 144);
peakEta_11_1_V <= s_INPUT_LINK_ARR( 3 )(156 downto 154);
peakPhi_11_1_V <= s_INPUT_LINK_ARR( 3 )(159 downto 157);
ClusterET_11_2_V <= s_INPUT_LINK_ARR( 3 )(169 downto 160);
peakEta_11_2_V <= s_INPUT_LINK_ARR( 3 )(172 downto 170);
peakPhi_11_2_V <= s_INPUT_LINK_ARR( 3 )(175 downto 173);
ClusterET_11_3_V <= s_INPUT_LINK_ARR( 3 )(185 downto 176);
peakEta_11_3_V <= s_INPUT_LINK_ARR( 3 )(188 downto 186);
peakPhi_11_3_V <= s_INPUT_LINK_ARR( 3 )(191 downto 189);
ClusterET_12_0_V <= s_INPUT_LINK_ARR( 4 )(9 downto 0);
peakEta_12_0_V <= s_INPUT_LINK_ARR( 4 )(12 downto 10);
peakPhi_12_0_V <= s_INPUT_LINK_ARR( 4 )(15 downto 13);
ClusterET_12_1_V <= s_INPUT_LINK_ARR( 4 )(25 downto 16);
peakEta_12_1_V <= s_INPUT_LINK_ARR( 4 )(28 downto 26);
peakPhi_12_1_V <= s_INPUT_LINK_ARR( 4 )(31 downto 29);
ClusterET_12_2_V <= s_INPUT_LINK_ARR( 4 )(41 downto 32);
peakEta_12_2_V <= s_INPUT_LINK_ARR( 4 )(44 downto 42);
peakPhi_12_2_V <= s_INPUT_LINK_ARR( 4 )(47 downto 45);
ClusterET_12_3_V <= s_INPUT_LINK_ARR( 4 )(57 downto 48);
peakEta_12_3_V <= s_INPUT_LINK_ARR( 4 )(60 downto 58);
peakPhi_12_3_V <= s_INPUT_LINK_ARR( 4 )(63 downto 61);
ClusterET_13_0_V <= s_INPUT_LINK_ARR( 4 )(73 downto 64);
peakEta_13_0_V <= s_INPUT_LINK_ARR( 4 )(76 downto 74);
peakPhi_13_0_V <= s_INPUT_LINK_ARR( 4 )(79 downto 77);
ClusterET_13_1_V <= s_INPUT_LINK_ARR( 4 )(89 downto 80);
peakEta_13_1_V <= s_INPUT_LINK_ARR( 4 )(92 downto 90);
peakPhi_13_1_V <= s_INPUT_LINK_ARR( 4 )(95 downto 93);
ClusterET_13_2_V <= s_INPUT_LINK_ARR( 4 )(105 downto 96);
peakEta_13_2_V <= s_INPUT_LINK_ARR( 4 )(108 downto 106);
peakPhi_13_2_V <= s_INPUT_LINK_ARR( 4 )(111 downto 109);
ClusterET_13_3_V <= s_INPUT_LINK_ARR( 4 )(121 downto 112);
peakEta_13_3_V <= s_INPUT_LINK_ARR( 4 )(124 downto 122);
peakPhi_13_3_V <= s_INPUT_LINK_ARR( 4 )(127 downto 125);
ClusterET_14_0_V <= s_INPUT_LINK_ARR( 4 )(137 downto 128);
peakEta_14_0_V <= s_INPUT_LINK_ARR( 4 )(140 downto 138);
peakPhi_14_0_V <= s_INPUT_LINK_ARR( 4 )(143 downto 141);
ClusterET_14_1_V <= s_INPUT_LINK_ARR( 4 )(153 downto 144);
peakEta_14_1_V <= s_INPUT_LINK_ARR( 4 )(156 downto 154);
peakPhi_14_1_V <= s_INPUT_LINK_ARR( 4 )(159 downto 157);
ClusterET_14_2_V <= s_INPUT_LINK_ARR( 4 )(169 downto 160);
peakEta_14_2_V <= s_INPUT_LINK_ARR( 4 )(172 downto 170);
peakPhi_14_2_V <= s_INPUT_LINK_ARR( 4 )(175 downto 173);
ClusterET_14_3_V <= s_INPUT_LINK_ARR( 4 )(185 downto 176);
peakEta_14_3_V <= s_INPUT_LINK_ARR( 4 )(188 downto 186);
peakPhi_14_3_V <= s_INPUT_LINK_ARR( 4 )(191 downto 189);
ClusterET_15_0_V <= s_INPUT_LINK_ARR( 5 )(9 downto 0);
peakEta_15_0_V <= s_INPUT_LINK_ARR( 5 )(12 downto 10);
peakPhi_15_0_V <= s_INPUT_LINK_ARR( 5 )(15 downto 13);
ClusterET_15_1_V <= s_INPUT_LINK_ARR( 5 )(25 downto 16);
peakEta_15_1_V <= s_INPUT_LINK_ARR( 5 )(28 downto 26);
peakPhi_15_1_V <= s_INPUT_LINK_ARR( 5 )(31 downto 29);
ClusterET_15_2_V <= s_INPUT_LINK_ARR( 5 )(41 downto 32);
peakEta_15_2_V <= s_INPUT_LINK_ARR( 5 )(44 downto 42);
peakPhi_15_2_V <= s_INPUT_LINK_ARR( 5 )(47 downto 45);
ClusterET_15_3_V <= s_INPUT_LINK_ARR( 5 )(57 downto 48);
peakEta_15_3_V <= s_INPUT_LINK_ARR( 5 )(60 downto 58);
peakPhi_15_3_V <= s_INPUT_LINK_ARR( 5 )(63 downto 61);
ClusterET_16_0_V <= s_INPUT_LINK_ARR( 5 )(73 downto 64);
peakEta_16_0_V <= s_INPUT_LINK_ARR( 5 )(76 downto 74);
peakPhi_16_0_V <= s_INPUT_LINK_ARR( 5 )(79 downto 77);
ClusterET_16_1_V <= s_INPUT_LINK_ARR( 5 )(89 downto 80);
peakEta_16_1_V <= s_INPUT_LINK_ARR( 5 )(92 downto 90);
peakPhi_16_1_V <= s_INPUT_LINK_ARR( 5 )(95 downto 93);
ClusterET_16_2_V <= s_INPUT_LINK_ARR( 5 )(105 downto 96);
peakEta_16_2_V <= s_INPUT_LINK_ARR( 5 )(108 downto 106);
peakPhi_16_2_V <= s_INPUT_LINK_ARR( 5 )(111 downto 109);
ClusterET_16_3_V <= s_INPUT_LINK_ARR( 5 )(121 downto 112);
peakEta_16_3_V <= s_INPUT_LINK_ARR( 5 )(124 downto 122);
peakPhi_16_3_V <= s_INPUT_LINK_ARR( 5 )(127 downto 125);


trackPT_0_V <= s_INPUT_LINK_ARR( 5 )(137 downto 128);
trackPT_1_V <= s_INPUT_LINK_ARR( 5 )(153 downto 144);
trackPT_2_V <= s_INPUT_LINK_ARR( 5 )(169 downto 160);
trackPT_3_V <= s_INPUT_LINK_ARR( 5 )(185 downto 176);
trackPT_4_V <= s_INPUT_LINK_ARR( 6 )(9 downto 0);
trackPT_5_V <= s_INPUT_LINK_ARR( 6 )(25 downto 16);
trackPT_6_V <= s_INPUT_LINK_ARR( 6 )(41 downto 32);
trackPT_7_V <= s_INPUT_LINK_ARR( 6 )(57 downto 48);
trackPT_8_V <= s_INPUT_LINK_ARR( 6 )(73 downto 64);
trackPT_9_V <= s_INPUT_LINK_ARR( 6 )(89 downto 80);


trackEta_0_V <= s_INPUT_LINK_ARR( 6 )(104 downto 96);
trackEta_1_V <= s_INPUT_LINK_ARR( 6 )(120 downto 112);
trackEta_2_V <= s_INPUT_LINK_ARR( 6 )(136 downto 128);
trackEta_3_V <= s_INPUT_LINK_ARR( 6 )(152 downto 144);
trackEta_4_V <= s_INPUT_LINK_ARR( 6 )(168 downto 160);
trackEta_5_V <= s_INPUT_LINK_ARR( 6 )(184 downto 176);
trackEta_6_V <= s_INPUT_LINK_ARR( 7 )(8 downto 0);
trackEta_7_V <= s_INPUT_LINK_ARR( 7 )(24 downto 16);
trackEta_8_V <= s_INPUT_LINK_ARR( 7 )(40 downto 32);
trackEta_9_V <= s_INPUT_LINK_ARR( 7 )(56 downto 48);


trackPhi_0_V <= s_INPUT_LINK_ARR( 7 )(73 downto 64);
trackPhi_1_V <= s_INPUT_LINK_ARR( 7 )(89 downto 80);
trackPhi_2_V <= s_INPUT_LINK_ARR( 7 )(105 downto 96);
trackPhi_3_V <= s_INPUT_LINK_ARR( 7 )(121 downto 112);
trackPhi_4_V <= s_INPUT_LINK_ARR( 7 )(137 downto 128);
trackPhi_5_V <= s_INPUT_LINK_ARR( 7 )(153 downto 144);
trackPhi_6_V <= s_INPUT_LINK_ARR( 7 )(169 downto 160);
trackPhi_7_V <= s_INPUT_LINK_ARR( 7 )(185 downto 176);
trackPhi_8_V <= s_INPUT_LINK_ARR( 8 )(9 downto 0);
trackPhi_9_V <= s_INPUT_LINK_ARR( 8 )(25 downto 16);


s_OUTPUT_LINK_ARR( 0 )(9 downto 0) <= output_linkedTrackPT_0_V ;
s_OUTPUT_LINK_ARR( 0 )(25 downto 16) <= output_linkedTrackPT_1_V ;
s_OUTPUT_LINK_ARR( 0 )(41 downto 32) <= output_linkedTrackPT_2_V ;
s_OUTPUT_LINK_ARR( 0 )(57 downto 48) <= output_linkedTrackPT_3_V ;
s_OUTPUT_LINK_ARR( 0 )(73 downto 64) <= output_linkedTrackPT_4_V ;
s_OUTPUT_LINK_ARR( 0 )(89 downto 80) <= output_linkedTrackPT_5_V ;
s_OUTPUT_LINK_ARR( 0 )(105 downto 96) <= output_linkedTrackPT_6_V ;
s_OUTPUT_LINK_ARR( 0 )(121 downto 112) <= output_linkedTrackPT_7_V ;
s_OUTPUT_LINK_ARR( 0 )(137 downto 128) <= output_linkedTrackPT_8_V ;
s_OUTPUT_LINK_ARR( 0 )(153 downto 144) <= output_linkedTrackPT_9_V ;


s_OUTPUT_LINK_ARR( 0 )(168 downto 160) <= output_linkedTrackEta_0_V ;
s_OUTPUT_LINK_ARR( 0 )(184 downto 176) <= output_linkedTrackEta_1_V ;
s_OUTPUT_LINK_ARR( 1 )(8 downto 0) <= output_linkedTrackEta_2_V ;
s_OUTPUT_LINK_ARR( 1 )(24 downto 16) <= output_linkedTrackEta_3_V ;
s_OUTPUT_LINK_ARR( 1 )(40 downto 32) <= output_linkedTrackEta_4_V ;
s_OUTPUT_LINK_ARR( 1 )(56 downto 48) <= output_linkedTrackEta_5_V ;
s_OUTPUT_LINK_ARR( 1 )(72 downto 64) <= output_linkedTrackEta_6_V ;
s_OUTPUT_LINK_ARR( 1 )(88 downto 80) <= output_linkedTrackEta_7_V ;
s_OUTPUT_LINK_ARR( 1 )(104 downto 96) <= output_linkedTrackEta_8_V ;
s_OUTPUT_LINK_ARR( 1 )(120 downto 112) <= output_linkedTrackEta_9_V ;


s_OUTPUT_LINK_ARR( 1 )(137 downto 128) <= output_linkedTrackPhi_0_V ;
s_OUTPUT_LINK_ARR( 1 )(153 downto 144) <= output_linkedTrackPhi_1_V ;
s_OUTPUT_LINK_ARR( 1 )(169 downto 160) <= output_linkedTrackPhi_2_V ;
s_OUTPUT_LINK_ARR( 1 )(185 downto 176) <= output_linkedTrackPhi_3_V ;
s_OUTPUT_LINK_ARR( 2 )(9 downto 0) <= output_linkedTrackPhi_4_V ;
s_OUTPUT_LINK_ARR( 2 )(25 downto 16) <= output_linkedTrackPhi_5_V ;
s_OUTPUT_LINK_ARR( 2 )(41 downto 32) <= output_linkedTrackPhi_6_V ;
s_OUTPUT_LINK_ARR( 2 )(57 downto 48) <= output_linkedTrackPhi_7_V ;
s_OUTPUT_LINK_ARR( 2 )(73 downto 64) <= output_linkedTrackPhi_8_V ;
s_OUTPUT_LINK_ARR( 2 )(89 downto 80) <= output_linkedTrackPhi_9_V ;


s_OUTPUT_LINK_ARR( 2 )(103 downto 96) <= output_linkedTrackQuality_0_V ;
s_OUTPUT_LINK_ARR( 2 )(119 downto 112) <= output_linkedTrackQuality_1_V ;
s_OUTPUT_LINK_ARR( 2 )(135 downto 128) <= output_linkedTrackQuality_2_V ;
s_OUTPUT_LINK_ARR( 2 )(151 downto 144) <= output_linkedTrackQuality_3_V ;
s_OUTPUT_LINK_ARR( 2 )(167 downto 160) <= output_linkedTrackQuality_4_V ;
s_OUTPUT_LINK_ARR( 2 )(183 downto 176) <= output_linkedTrackQuality_5_V ;
s_OUTPUT_LINK_ARR( 3 )(7 downto 0) <= output_linkedTrackQuality_6_V ;
s_OUTPUT_LINK_ARR( 3 )(23 downto 16) <= output_linkedTrackQuality_7_V ;
s_OUTPUT_LINK_ARR( 3 )(39 downto 32) <= output_linkedTrackQuality_8_V ;
s_OUTPUT_LINK_ARR( 3 )(55 downto 48) <= output_linkedTrackQuality_9_V ;


s_OUTPUT_LINK_ARR( 3 )(73 downto 64) <= output_neutralClusterET_0_V ;
s_OUTPUT_LINK_ARR( 3 )(89 downto 80) <= output_neutralClusterET_1_V ;
s_OUTPUT_LINK_ARR( 3 )(105 downto 96) <= output_neutralClusterET_2_V ;
s_OUTPUT_LINK_ARR( 3 )(121 downto 112) <= output_neutralClusterET_3_V ;
s_OUTPUT_LINK_ARR( 3 )(137 downto 128) <= output_neutralClusterET_4_V ;
s_OUTPUT_LINK_ARR( 3 )(153 downto 144) <= output_neutralClusterET_5_V ;
s_OUTPUT_LINK_ARR( 3 )(169 downto 160) <= output_neutralClusterET_6_V ;
s_OUTPUT_LINK_ARR( 3 )(185 downto 176) <= output_neutralClusterET_7_V ;
s_OUTPUT_LINK_ARR( 4 )(9 downto 0) <= output_neutralClusterET_8_V ;
s_OUTPUT_LINK_ARR( 4 )(25 downto 16) <= output_neutralClusterET_9_V ;
s_OUTPUT_LINK_ARR( 4 )(41 downto 32) <= output_neutralClusterET_10_V ;
s_OUTPUT_LINK_ARR( 4 )(57 downto 48) <= output_neutralClusterET_11_V ;
s_OUTPUT_LINK_ARR( 4 )(73 downto 64) <= output_neutralClusterET_12_V ;
s_OUTPUT_LINK_ARR( 4 )(89 downto 80) <= output_neutralClusterET_13_V ;
s_OUTPUT_LINK_ARR( 4 )(105 downto 96) <= output_neutralClusterET_14_V ;
s_OUTPUT_LINK_ARR( 4 )(121 downto 112) <= output_neutralClusterET_15_V ;
s_OUTPUT_LINK_ARR( 4 )(137 downto 128) <= output_neutralClusterET_16_V ;
s_OUTPUT_LINK_ARR( 4 )(153 downto 144) <= output_neutralClusterET_17_V ;
s_OUTPUT_LINK_ARR( 4 )(169 downto 160) <= output_neutralClusterET_18_V ;
s_OUTPUT_LINK_ARR( 4 )(185 downto 176) <= output_neutralClusterET_19_V ;
s_OUTPUT_LINK_ARR( 5 )(9 downto 0) <= output_neutralClusterET_20_V ;
s_OUTPUT_LINK_ARR( 5 )(25 downto 16) <= output_neutralClusterET_21_V ;
s_OUTPUT_LINK_ARR( 5 )(41 downto 32) <= output_neutralClusterET_22_V ;
s_OUTPUT_LINK_ARR( 5 )(57 downto 48) <= output_neutralClusterET_23_V ;
s_OUTPUT_LINK_ARR( 5 )(73 downto 64) <= output_neutralClusterET_24_V ;
s_OUTPUT_LINK_ARR( 5 )(89 downto 80) <= output_neutralClusterET_25_V ;
s_OUTPUT_LINK_ARR( 5 )(105 downto 96) <= output_neutralClusterET_26_V ;
s_OUTPUT_LINK_ARR( 5 )(121 downto 112) <= output_neutralClusterET_27_V ;
s_OUTPUT_LINK_ARR( 5 )(137 downto 128) <= output_neutralClusterET_28_V ;
s_OUTPUT_LINK_ARR( 5 )(153 downto 144) <= output_neutralClusterET_29_V ;
s_OUTPUT_LINK_ARR( 5 )(169 downto 160) <= output_neutralClusterET_30_V ;
s_OUTPUT_LINK_ARR( 5 )(185 downto 176) <= output_neutralClusterET_31_V ;
s_OUTPUT_LINK_ARR( 6 )(9 downto 0) <= output_neutralClusterET_32_V ;
s_OUTPUT_LINK_ARR( 6 )(25 downto 16) <= output_neutralClusterET_33_V ;
s_OUTPUT_LINK_ARR( 6 )(41 downto 32) <= output_neutralClusterET_34_V ;
s_OUTPUT_LINK_ARR( 6 )(57 downto 48) <= output_neutralClusterET_35_V ;
s_OUTPUT_LINK_ARR( 6 )(73 downto 64) <= output_neutralClusterET_36_V ;
s_OUTPUT_LINK_ARR( 6 )(89 downto 80) <= output_neutralClusterET_37_V ;
s_OUTPUT_LINK_ARR( 6 )(105 downto 96) <= output_neutralClusterET_38_V ;
s_OUTPUT_LINK_ARR( 6 )(121 downto 112) <= output_neutralClusterET_39_V ;
s_OUTPUT_LINK_ARR( 6 )(137 downto 128) <= output_neutralClusterET_40_V ;
s_OUTPUT_LINK_ARR( 6 )(153 downto 144) <= output_neutralClusterET_41_V ;
s_OUTPUT_LINK_ARR( 6 )(169 downto 160) <= output_neutralClusterET_42_V ;
s_OUTPUT_LINK_ARR( 6 )(185 downto 176) <= output_neutralClusterET_43_V ;
s_OUTPUT_LINK_ARR( 7 )(9 downto 0) <= output_neutralClusterET_44_V ;
s_OUTPUT_LINK_ARR( 7 )(25 downto 16) <= output_neutralClusterET_45_V ;
s_OUTPUT_LINK_ARR( 7 )(41 downto 32) <= output_neutralClusterET_46_V ;
s_OUTPUT_LINK_ARR( 7 )(57 downto 48) <= output_neutralClusterET_47_V ;
s_OUTPUT_LINK_ARR( 7 )(73 downto 64) <= output_neutralClusterET_48_V ;
s_OUTPUT_LINK_ARR( 7 )(89 downto 80) <= output_neutralClusterET_49_V ;
s_OUTPUT_LINK_ARR( 7 )(105 downto 96) <= output_neutralClusterET_50_V ;
s_OUTPUT_LINK_ARR( 7 )(121 downto 112) <= output_neutralClusterET_51_V ;
s_OUTPUT_LINK_ARR( 7 )(137 downto 128) <= output_neutralClusterET_52_V ;
s_OUTPUT_LINK_ARR( 7 )(153 downto 144) <= output_neutralClusterET_53_V ;
s_OUTPUT_LINK_ARR( 7 )(169 downto 160) <= output_neutralClusterET_54_V ;
s_OUTPUT_LINK_ARR( 7 )(185 downto 176) <= output_neutralClusterET_55_V ;
s_OUTPUT_LINK_ARR( 8 )(9 downto 0) <= output_neutralClusterET_56_V ;
s_OUTPUT_LINK_ARR( 8 )(25 downto 16) <= output_neutralClusterET_57_V ;
s_OUTPUT_LINK_ARR( 8 )(41 downto 32) <= output_neutralClusterET_58_V ;
s_OUTPUT_LINK_ARR( 8 )(57 downto 48) <= output_neutralClusterET_59_V ;
s_OUTPUT_LINK_ARR( 8 )(73 downto 64) <= output_neutralClusterET_60_V ;
s_OUTPUT_LINK_ARR( 8 )(89 downto 80) <= output_neutralClusterET_61_V ;
s_OUTPUT_LINK_ARR( 8 )(105 downto 96) <= output_neutralClusterET_62_V ;
s_OUTPUT_LINK_ARR( 8 )(121 downto 112) <= output_neutralClusterET_63_V ;
s_OUTPUT_LINK_ARR( 8 )(137 downto 128) <= output_neutralClusterET_64_V ;
s_OUTPUT_LINK_ARR( 8 )(153 downto 144) <= output_neutralClusterET_65_V ;
s_OUTPUT_LINK_ARR( 8 )(169 downto 160) <= output_neutralClusterET_66_V ;
s_OUTPUT_LINK_ARR( 8 )(185 downto 176) <= output_neutralClusterET_67_V ;


s_OUTPUT_LINK_ARR( 9 )(8 downto 0) <= output_neutralClusterEta_0_V ;
s_OUTPUT_LINK_ARR( 9 )(24 downto 16) <= output_neutralClusterEta_1_V ;
s_OUTPUT_LINK_ARR( 9 )(40 downto 32) <= output_neutralClusterEta_2_V ;
s_OUTPUT_LINK_ARR( 9 )(56 downto 48) <= output_neutralClusterEta_3_V ;
s_OUTPUT_LINK_ARR( 9 )(72 downto 64) <= output_neutralClusterEta_4_V ;
s_OUTPUT_LINK_ARR( 9 )(88 downto 80) <= output_neutralClusterEta_5_V ;
s_OUTPUT_LINK_ARR( 9 )(104 downto 96) <= output_neutralClusterEta_6_V ;
s_OUTPUT_LINK_ARR( 9 )(120 downto 112) <= output_neutralClusterEta_7_V ;
s_OUTPUT_LINK_ARR( 9 )(136 downto 128) <= output_neutralClusterEta_8_V ;
s_OUTPUT_LINK_ARR( 9 )(152 downto 144) <= output_neutralClusterEta_9_V ;
s_OUTPUT_LINK_ARR( 9 )(168 downto 160) <= output_neutralClusterEta_10_V ;
s_OUTPUT_LINK_ARR( 9 )(184 downto 176) <= output_neutralClusterEta_11_V ;
s_OUTPUT_LINK_ARR( 10 )(8 downto 0) <= output_neutralClusterEta_12_V ;
s_OUTPUT_LINK_ARR( 10 )(24 downto 16) <= output_neutralClusterEta_13_V ;
s_OUTPUT_LINK_ARR( 10 )(40 downto 32) <= output_neutralClusterEta_14_V ;
s_OUTPUT_LINK_ARR( 10 )(56 downto 48) <= output_neutralClusterEta_15_V ;
s_OUTPUT_LINK_ARR( 10 )(72 downto 64) <= output_neutralClusterEta_16_V ;
s_OUTPUT_LINK_ARR( 10 )(88 downto 80) <= output_neutralClusterEta_17_V ;
s_OUTPUT_LINK_ARR( 10 )(104 downto 96) <= output_neutralClusterEta_18_V ;
s_OUTPUT_LINK_ARR( 10 )(120 downto 112) <= output_neutralClusterEta_19_V ;
s_OUTPUT_LINK_ARR( 10 )(136 downto 128) <= output_neutralClusterEta_20_V ;
s_OUTPUT_LINK_ARR( 10 )(152 downto 144) <= output_neutralClusterEta_21_V ;
s_OUTPUT_LINK_ARR( 10 )(168 downto 160) <= output_neutralClusterEta_22_V ;
s_OUTPUT_LINK_ARR( 10 )(184 downto 176) <= output_neutralClusterEta_23_V ;
s_OUTPUT_LINK_ARR( 11 )(8 downto 0) <= output_neutralClusterEta_24_V ;
s_OUTPUT_LINK_ARR( 11 )(24 downto 16) <= output_neutralClusterEta_25_V ;
s_OUTPUT_LINK_ARR( 11 )(40 downto 32) <= output_neutralClusterEta_26_V ;
s_OUTPUT_LINK_ARR( 11 )(56 downto 48) <= output_neutralClusterEta_27_V ;
s_OUTPUT_LINK_ARR( 11 )(72 downto 64) <= output_neutralClusterEta_28_V ;
s_OUTPUT_LINK_ARR( 11 )(88 downto 80) <= output_neutralClusterEta_29_V ;
s_OUTPUT_LINK_ARR( 11 )(104 downto 96) <= output_neutralClusterEta_30_V ;
s_OUTPUT_LINK_ARR( 11 )(120 downto 112) <= output_neutralClusterEta_31_V ;
s_OUTPUT_LINK_ARR( 11 )(136 downto 128) <= output_neutralClusterEta_32_V ;
s_OUTPUT_LINK_ARR( 11 )(152 downto 144) <= output_neutralClusterEta_33_V ;
s_OUTPUT_LINK_ARR( 11 )(168 downto 160) <= output_neutralClusterEta_34_V ;
s_OUTPUT_LINK_ARR( 11 )(184 downto 176) <= output_neutralClusterEta_35_V ;
s_OUTPUT_LINK_ARR( 12 )(8 downto 0) <= output_neutralClusterEta_36_V ;
s_OUTPUT_LINK_ARR( 12 )(24 downto 16) <= output_neutralClusterEta_37_V ;
s_OUTPUT_LINK_ARR( 12 )(40 downto 32) <= output_neutralClusterEta_38_V ;
s_OUTPUT_LINK_ARR( 12 )(56 downto 48) <= output_neutralClusterEta_39_V ;
s_OUTPUT_LINK_ARR( 12 )(72 downto 64) <= output_neutralClusterEta_40_V ;
s_OUTPUT_LINK_ARR( 12 )(88 downto 80) <= output_neutralClusterEta_41_V ;
s_OUTPUT_LINK_ARR( 12 )(104 downto 96) <= output_neutralClusterEta_42_V ;
s_OUTPUT_LINK_ARR( 12 )(120 downto 112) <= output_neutralClusterEta_43_V ;
s_OUTPUT_LINK_ARR( 12 )(136 downto 128) <= output_neutralClusterEta_44_V ;
s_OUTPUT_LINK_ARR( 12 )(152 downto 144) <= output_neutralClusterEta_45_V ;
s_OUTPUT_LINK_ARR( 12 )(168 downto 160) <= output_neutralClusterEta_46_V ;
s_OUTPUT_LINK_ARR( 12 )(184 downto 176) <= output_neutralClusterEta_47_V ;
s_OUTPUT_LINK_ARR( 13 )(8 downto 0) <= output_neutralClusterEta_48_V ;
s_OUTPUT_LINK_ARR( 13 )(24 downto 16) <= output_neutralClusterEta_49_V ;
s_OUTPUT_LINK_ARR( 13 )(40 downto 32) <= output_neutralClusterEta_50_V ;
s_OUTPUT_LINK_ARR( 13 )(56 downto 48) <= output_neutralClusterEta_51_V ;
s_OUTPUT_LINK_ARR( 13 )(72 downto 64) <= output_neutralClusterEta_52_V ;
s_OUTPUT_LINK_ARR( 13 )(88 downto 80) <= output_neutralClusterEta_53_V ;
s_OUTPUT_LINK_ARR( 13 )(104 downto 96) <= output_neutralClusterEta_54_V ;
s_OUTPUT_LINK_ARR( 13 )(120 downto 112) <= output_neutralClusterEta_55_V ;
s_OUTPUT_LINK_ARR( 13 )(136 downto 128) <= output_neutralClusterEta_56_V ;
s_OUTPUT_LINK_ARR( 13 )(152 downto 144) <= output_neutralClusterEta_57_V ;
s_OUTPUT_LINK_ARR( 13 )(168 downto 160) <= output_neutralClusterEta_58_V ;
s_OUTPUT_LINK_ARR( 13 )(184 downto 176) <= output_neutralClusterEta_59_V ;
s_OUTPUT_LINK_ARR( 14 )(8 downto 0) <= output_neutralClusterEta_60_V ;
s_OUTPUT_LINK_ARR( 14 )(24 downto 16) <= output_neutralClusterEta_61_V ;
s_OUTPUT_LINK_ARR( 14 )(40 downto 32) <= output_neutralClusterEta_62_V ;
s_OUTPUT_LINK_ARR( 14 )(56 downto 48) <= output_neutralClusterEta_63_V ;
s_OUTPUT_LINK_ARR( 14 )(72 downto 64) <= output_neutralClusterEta_64_V ;
s_OUTPUT_LINK_ARR( 14 )(88 downto 80) <= output_neutralClusterEta_65_V ;
s_OUTPUT_LINK_ARR( 14 )(104 downto 96) <= output_neutralClusterEta_66_V ;
s_OUTPUT_LINK_ARR( 14 )(120 downto 112) <= output_neutralClusterEta_67_V ;


s_OUTPUT_LINK_ARR( 14 )(137 downto 128) <= output_neutralClusterPhi_0_V ;
s_OUTPUT_LINK_ARR( 14 )(153 downto 144) <= output_neutralClusterPhi_1_V ;
s_OUTPUT_LINK_ARR( 14 )(169 downto 160) <= output_neutralClusterPhi_2_V ;
s_OUTPUT_LINK_ARR( 14 )(185 downto 176) <= output_neutralClusterPhi_3_V ;
s_OUTPUT_LINK_ARR( 15 )(9 downto 0) <= output_neutralClusterPhi_4_V ;
s_OUTPUT_LINK_ARR( 15 )(25 downto 16) <= output_neutralClusterPhi_5_V ;
s_OUTPUT_LINK_ARR( 15 )(41 downto 32) <= output_neutralClusterPhi_6_V ;
s_OUTPUT_LINK_ARR( 15 )(57 downto 48) <= output_neutralClusterPhi_7_V ;
s_OUTPUT_LINK_ARR( 15 )(73 downto 64) <= output_neutralClusterPhi_8_V ;
s_OUTPUT_LINK_ARR( 15 )(89 downto 80) <= output_neutralClusterPhi_9_V ;
s_OUTPUT_LINK_ARR( 15 )(105 downto 96) <= output_neutralClusterPhi_10_V ;
s_OUTPUT_LINK_ARR( 15 )(121 downto 112) <= output_neutralClusterPhi_11_V ;
s_OUTPUT_LINK_ARR( 15 )(137 downto 128) <= output_neutralClusterPhi_12_V ;
s_OUTPUT_LINK_ARR( 15 )(153 downto 144) <= output_neutralClusterPhi_13_V ;
s_OUTPUT_LINK_ARR( 15 )(169 downto 160) <= output_neutralClusterPhi_14_V ;
s_OUTPUT_LINK_ARR( 15 )(185 downto 176) <= output_neutralClusterPhi_15_V ;
s_OUTPUT_LINK_ARR( 16 )(9 downto 0) <= output_neutralClusterPhi_16_V ;
s_OUTPUT_LINK_ARR( 16 )(25 downto 16) <= output_neutralClusterPhi_17_V ;
s_OUTPUT_LINK_ARR( 16 )(41 downto 32) <= output_neutralClusterPhi_18_V ;
s_OUTPUT_LINK_ARR( 16 )(57 downto 48) <= output_neutralClusterPhi_19_V ;
s_OUTPUT_LINK_ARR( 16 )(73 downto 64) <= output_neutralClusterPhi_20_V ;
s_OUTPUT_LINK_ARR( 16 )(89 downto 80) <= output_neutralClusterPhi_21_V ;
s_OUTPUT_LINK_ARR( 16 )(105 downto 96) <= output_neutralClusterPhi_22_V ;
s_OUTPUT_LINK_ARR( 16 )(121 downto 112) <= output_neutralClusterPhi_23_V ;
s_OUTPUT_LINK_ARR( 16 )(137 downto 128) <= output_neutralClusterPhi_24_V ;
s_OUTPUT_LINK_ARR( 16 )(153 downto 144) <= output_neutralClusterPhi_25_V ;
s_OUTPUT_LINK_ARR( 16 )(169 downto 160) <= output_neutralClusterPhi_26_V ;
s_OUTPUT_LINK_ARR( 16 )(185 downto 176) <= output_neutralClusterPhi_27_V ;
s_OUTPUT_LINK_ARR( 17 )(9 downto 0) <= output_neutralClusterPhi_28_V ;
s_OUTPUT_LINK_ARR( 17 )(25 downto 16) <= output_neutralClusterPhi_29_V ;
s_OUTPUT_LINK_ARR( 17 )(41 downto 32) <= output_neutralClusterPhi_30_V ;
s_OUTPUT_LINK_ARR( 17 )(57 downto 48) <= output_neutralClusterPhi_31_V ;
s_OUTPUT_LINK_ARR( 17 )(73 downto 64) <= output_neutralClusterPhi_32_V ;
s_OUTPUT_LINK_ARR( 17 )(89 downto 80) <= output_neutralClusterPhi_33_V ;
s_OUTPUT_LINK_ARR( 17 )(105 downto 96) <= output_neutralClusterPhi_34_V ;
s_OUTPUT_LINK_ARR( 17 )(121 downto 112) <= output_neutralClusterPhi_35_V ;
s_OUTPUT_LINK_ARR( 17 )(137 downto 128) <= output_neutralClusterPhi_36_V ;
s_OUTPUT_LINK_ARR( 17 )(153 downto 144) <= output_neutralClusterPhi_37_V ;
s_OUTPUT_LINK_ARR( 17 )(169 downto 160) <= output_neutralClusterPhi_38_V ;
s_OUTPUT_LINK_ARR( 17 )(185 downto 176) <= output_neutralClusterPhi_39_V ;
s_OUTPUT_LINK_ARR( 18 )(9 downto 0) <= output_neutralClusterPhi_40_V ;
s_OUTPUT_LINK_ARR( 18 )(25 downto 16) <= output_neutralClusterPhi_41_V ;
s_OUTPUT_LINK_ARR( 18 )(41 downto 32) <= output_neutralClusterPhi_42_V ;
s_OUTPUT_LINK_ARR( 18 )(57 downto 48) <= output_neutralClusterPhi_43_V ;
s_OUTPUT_LINK_ARR( 18 )(73 downto 64) <= output_neutralClusterPhi_44_V ;
s_OUTPUT_LINK_ARR( 18 )(89 downto 80) <= output_neutralClusterPhi_45_V ;
s_OUTPUT_LINK_ARR( 18 )(105 downto 96) <= output_neutralClusterPhi_46_V ;
s_OUTPUT_LINK_ARR( 18 )(121 downto 112) <= output_neutralClusterPhi_47_V ;
s_OUTPUT_LINK_ARR( 18 )(137 downto 128) <= output_neutralClusterPhi_48_V ;
s_OUTPUT_LINK_ARR( 18 )(153 downto 144) <= output_neutralClusterPhi_49_V ;
s_OUTPUT_LINK_ARR( 18 )(169 downto 160) <= output_neutralClusterPhi_50_V ;
s_OUTPUT_LINK_ARR( 18 )(185 downto 176) <= output_neutralClusterPhi_51_V ;
s_OUTPUT_LINK_ARR( 19 )(9 downto 0) <= output_neutralClusterPhi_52_V ;
s_OUTPUT_LINK_ARR( 19 )(25 downto 16) <= output_neutralClusterPhi_53_V ;
s_OUTPUT_LINK_ARR( 19 )(41 downto 32) <= output_neutralClusterPhi_54_V ;
s_OUTPUT_LINK_ARR( 19 )(57 downto 48) <= output_neutralClusterPhi_55_V ;
s_OUTPUT_LINK_ARR( 19 )(73 downto 64) <= output_neutralClusterPhi_56_V ;
s_OUTPUT_LINK_ARR( 19 )(89 downto 80) <= output_neutralClusterPhi_57_V ;
s_OUTPUT_LINK_ARR( 19 )(105 downto 96) <= output_neutralClusterPhi_58_V ;
s_OUTPUT_LINK_ARR( 19 )(121 downto 112) <= output_neutralClusterPhi_59_V ;
s_OUTPUT_LINK_ARR( 19 )(137 downto 128) <= output_neutralClusterPhi_60_V ;
s_OUTPUT_LINK_ARR( 19 )(153 downto 144) <= output_neutralClusterPhi_61_V ;
s_OUTPUT_LINK_ARR( 19 )(169 downto 160) <= output_neutralClusterPhi_62_V ;
s_OUTPUT_LINK_ARR( 19 )(185 downto 176) <= output_neutralClusterPhi_63_V ;
s_OUTPUT_LINK_ARR( 20 )(9 downto 0) <= output_neutralClusterPhi_64_V ;
s_OUTPUT_LINK_ARR( 20 )(25 downto 16) <= output_neutralClusterPhi_65_V ;
s_OUTPUT_LINK_ARR( 20 )(41 downto 32) <= output_neutralClusterPhi_66_V ;
s_OUTPUT_LINK_ARR( 20 )(57 downto 48) <= output_neutralClusterPhi_67_V ;




------

-----------------------------------------------------------------------------
-- End User_Code
-----------------------------------------------------------------------------

end ctp7_top_arch;
